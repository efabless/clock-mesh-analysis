magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1260 -1260 1261 1261
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 1449762
string GDS_START 1449310
<< end >>

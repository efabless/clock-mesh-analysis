magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1288 -1260 1936 1357
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_2
timestamp 1633016201
transform 1 0 472 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_1
timestamp 1633016201
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_0
timestamp 1633016201
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_1
timestamp 1633016201
transform 1 0 648 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1633016201
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 676 97 676 97 0 FreeSans 300 0 0 0 S
flabel comment s 500 97 500 97 0 FreeSans 300 0 0 0 D
flabel comment s 324 97 324 97 0 FreeSans 300 0 0 0 S
flabel comment s 148 97 148 97 0 FreeSans 300 0 0 0 D
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 39944018
string GDS_START 39941218
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -2178 -1679 2412 16012
<< dnwell >>
rect -122 -335 1072 4993
<< nwell >>
rect -918 13930 952 14752
rect -918 5076 86 13930
rect -918 4908 1152 5076
rect -918 168 168 4908
rect 782 168 1152 4908
rect -918 -202 1152 168
rect -918 -419 964 -202
<< pwell >>
rect 228 228 722 4848
<< mvnmos >>
rect 415 3714 535 4714
rect 415 2593 535 3593
rect 415 1472 535 2472
rect 415 362 535 1362
<< mvndiff >>
rect 362 4702 415 4714
rect 362 4668 370 4702
rect 404 4668 415 4702
rect 362 4634 415 4668
rect 362 4600 370 4634
rect 404 4600 415 4634
rect 362 4566 415 4600
rect 362 4532 370 4566
rect 404 4532 415 4566
rect 362 4498 415 4532
rect 362 4464 370 4498
rect 404 4464 415 4498
rect 362 4430 415 4464
rect 362 4396 370 4430
rect 404 4396 415 4430
rect 362 4362 415 4396
rect 362 4328 370 4362
rect 404 4328 415 4362
rect 362 4294 415 4328
rect 362 4260 370 4294
rect 404 4260 415 4294
rect 362 4226 415 4260
rect 362 4192 370 4226
rect 404 4192 415 4226
rect 362 4158 415 4192
rect 362 4124 370 4158
rect 404 4124 415 4158
rect 362 4090 415 4124
rect 362 4056 370 4090
rect 404 4056 415 4090
rect 362 4022 415 4056
rect 362 3988 370 4022
rect 404 3988 415 4022
rect 362 3954 415 3988
rect 362 3920 370 3954
rect 404 3920 415 3954
rect 362 3886 415 3920
rect 362 3852 370 3886
rect 404 3852 415 3886
rect 362 3818 415 3852
rect 362 3784 370 3818
rect 404 3784 415 3818
rect 362 3714 415 3784
rect 535 4702 588 4714
rect 535 4668 546 4702
rect 580 4668 588 4702
rect 535 4634 588 4668
rect 535 4600 546 4634
rect 580 4600 588 4634
rect 535 4566 588 4600
rect 535 4532 546 4566
rect 580 4532 588 4566
rect 535 4498 588 4532
rect 535 4464 546 4498
rect 580 4464 588 4498
rect 535 4430 588 4464
rect 535 4396 546 4430
rect 580 4396 588 4430
rect 535 4362 588 4396
rect 535 4328 546 4362
rect 580 4328 588 4362
rect 535 4294 588 4328
rect 535 4260 546 4294
rect 580 4260 588 4294
rect 535 4226 588 4260
rect 535 4192 546 4226
rect 580 4192 588 4226
rect 535 4158 588 4192
rect 535 4124 546 4158
rect 580 4124 588 4158
rect 535 4090 588 4124
rect 535 4056 546 4090
rect 580 4056 588 4090
rect 535 4022 588 4056
rect 535 3988 546 4022
rect 580 3988 588 4022
rect 535 3954 588 3988
rect 535 3920 546 3954
rect 580 3920 588 3954
rect 535 3886 588 3920
rect 535 3852 546 3886
rect 580 3852 588 3886
rect 535 3818 588 3852
rect 535 3784 546 3818
rect 580 3784 588 3818
rect 535 3714 588 3784
rect 362 3581 415 3593
rect 362 3547 370 3581
rect 404 3547 415 3581
rect 362 3513 415 3547
rect 362 3479 370 3513
rect 404 3479 415 3513
rect 362 3445 415 3479
rect 362 3411 370 3445
rect 404 3411 415 3445
rect 362 3377 415 3411
rect 362 3343 370 3377
rect 404 3343 415 3377
rect 362 3309 415 3343
rect 362 3275 370 3309
rect 404 3275 415 3309
rect 362 3241 415 3275
rect 362 3207 370 3241
rect 404 3207 415 3241
rect 362 3173 415 3207
rect 362 3139 370 3173
rect 404 3139 415 3173
rect 362 3105 415 3139
rect 362 3071 370 3105
rect 404 3071 415 3105
rect 362 3037 415 3071
rect 362 3003 370 3037
rect 404 3003 415 3037
rect 362 2969 415 3003
rect 362 2935 370 2969
rect 404 2935 415 2969
rect 362 2901 415 2935
rect 362 2867 370 2901
rect 404 2867 415 2901
rect 362 2833 415 2867
rect 362 2799 370 2833
rect 404 2799 415 2833
rect 362 2765 415 2799
rect 362 2731 370 2765
rect 404 2731 415 2765
rect 362 2697 415 2731
rect 362 2663 370 2697
rect 404 2663 415 2697
rect 362 2593 415 2663
rect 535 3581 588 3593
rect 535 3547 546 3581
rect 580 3547 588 3581
rect 535 3513 588 3547
rect 535 3479 546 3513
rect 580 3479 588 3513
rect 535 3445 588 3479
rect 535 3411 546 3445
rect 580 3411 588 3445
rect 535 3377 588 3411
rect 535 3343 546 3377
rect 580 3343 588 3377
rect 535 3309 588 3343
rect 535 3275 546 3309
rect 580 3275 588 3309
rect 535 3241 588 3275
rect 535 3207 546 3241
rect 580 3207 588 3241
rect 535 3173 588 3207
rect 535 3139 546 3173
rect 580 3139 588 3173
rect 535 3105 588 3139
rect 535 3071 546 3105
rect 580 3071 588 3105
rect 535 3037 588 3071
rect 535 3003 546 3037
rect 580 3003 588 3037
rect 535 2969 588 3003
rect 535 2935 546 2969
rect 580 2935 588 2969
rect 535 2901 588 2935
rect 535 2867 546 2901
rect 580 2867 588 2901
rect 535 2833 588 2867
rect 535 2799 546 2833
rect 580 2799 588 2833
rect 535 2765 588 2799
rect 535 2731 546 2765
rect 580 2731 588 2765
rect 535 2697 588 2731
rect 535 2663 546 2697
rect 580 2663 588 2697
rect 535 2593 588 2663
rect 362 2460 415 2472
rect 362 2426 370 2460
rect 404 2426 415 2460
rect 362 2392 415 2426
rect 362 2358 370 2392
rect 404 2358 415 2392
rect 362 2324 415 2358
rect 362 2290 370 2324
rect 404 2290 415 2324
rect 362 2256 415 2290
rect 362 2222 370 2256
rect 404 2222 415 2256
rect 362 2188 415 2222
rect 362 2154 370 2188
rect 404 2154 415 2188
rect 362 2120 415 2154
rect 362 2086 370 2120
rect 404 2086 415 2120
rect 362 2052 415 2086
rect 362 2018 370 2052
rect 404 2018 415 2052
rect 362 1984 415 2018
rect 362 1950 370 1984
rect 404 1950 415 1984
rect 362 1916 415 1950
rect 362 1882 370 1916
rect 404 1882 415 1916
rect 362 1848 415 1882
rect 362 1814 370 1848
rect 404 1814 415 1848
rect 362 1780 415 1814
rect 362 1746 370 1780
rect 404 1746 415 1780
rect 362 1712 415 1746
rect 362 1678 370 1712
rect 404 1678 415 1712
rect 362 1644 415 1678
rect 362 1610 370 1644
rect 404 1610 415 1644
rect 362 1576 415 1610
rect 362 1542 370 1576
rect 404 1542 415 1576
rect 362 1472 415 1542
rect 535 2460 588 2472
rect 535 2426 546 2460
rect 580 2426 588 2460
rect 535 2392 588 2426
rect 535 2358 546 2392
rect 580 2358 588 2392
rect 535 2324 588 2358
rect 535 2290 546 2324
rect 580 2290 588 2324
rect 535 2256 588 2290
rect 535 2222 546 2256
rect 580 2222 588 2256
rect 535 2188 588 2222
rect 535 2154 546 2188
rect 580 2154 588 2188
rect 535 2120 588 2154
rect 535 2086 546 2120
rect 580 2086 588 2120
rect 535 2052 588 2086
rect 535 2018 546 2052
rect 580 2018 588 2052
rect 535 1984 588 2018
rect 535 1950 546 1984
rect 580 1950 588 1984
rect 535 1916 588 1950
rect 535 1882 546 1916
rect 580 1882 588 1916
rect 535 1848 588 1882
rect 535 1814 546 1848
rect 580 1814 588 1848
rect 535 1780 588 1814
rect 535 1746 546 1780
rect 580 1746 588 1780
rect 535 1712 588 1746
rect 535 1678 546 1712
rect 580 1678 588 1712
rect 535 1644 588 1678
rect 535 1610 546 1644
rect 580 1610 588 1644
rect 535 1576 588 1610
rect 535 1542 546 1576
rect 580 1542 588 1576
rect 535 1472 588 1542
rect 362 1292 415 1362
rect 362 1258 370 1292
rect 404 1258 415 1292
rect 362 1224 415 1258
rect 362 1190 370 1224
rect 404 1190 415 1224
rect 362 1156 415 1190
rect 362 1122 370 1156
rect 404 1122 415 1156
rect 362 1088 415 1122
rect 362 1054 370 1088
rect 404 1054 415 1088
rect 362 1020 415 1054
rect 362 986 370 1020
rect 404 986 415 1020
rect 362 952 415 986
rect 362 918 370 952
rect 404 918 415 952
rect 362 884 415 918
rect 362 850 370 884
rect 404 850 415 884
rect 362 816 415 850
rect 362 782 370 816
rect 404 782 415 816
rect 362 748 415 782
rect 362 714 370 748
rect 404 714 415 748
rect 362 680 415 714
rect 362 646 370 680
rect 404 646 415 680
rect 362 612 415 646
rect 362 578 370 612
rect 404 578 415 612
rect 362 544 415 578
rect 362 510 370 544
rect 404 510 415 544
rect 362 476 415 510
rect 362 442 370 476
rect 404 442 415 476
rect 362 408 415 442
rect 362 374 370 408
rect 404 374 415 408
rect 362 362 415 374
rect 535 1292 588 1362
rect 535 1258 546 1292
rect 580 1258 588 1292
rect 535 1224 588 1258
rect 535 1190 546 1224
rect 580 1190 588 1224
rect 535 1156 588 1190
rect 535 1122 546 1156
rect 580 1122 588 1156
rect 535 1088 588 1122
rect 535 1054 546 1088
rect 580 1054 588 1088
rect 535 1020 588 1054
rect 535 986 546 1020
rect 580 986 588 1020
rect 535 952 588 986
rect 535 918 546 952
rect 580 918 588 952
rect 535 884 588 918
rect 535 850 546 884
rect 580 850 588 884
rect 535 816 588 850
rect 535 782 546 816
rect 580 782 588 816
rect 535 748 588 782
rect 535 714 546 748
rect 580 714 588 748
rect 535 680 588 714
rect 535 646 546 680
rect 580 646 588 680
rect 535 612 588 646
rect 535 578 546 612
rect 580 578 588 612
rect 535 544 588 578
rect 535 510 546 544
rect 580 510 588 544
rect 535 476 588 510
rect 535 442 546 476
rect 580 442 588 476
rect 535 408 588 442
rect 535 374 546 408
rect 580 374 588 408
rect 535 362 588 374
<< mvndiffc >>
rect 370 4668 404 4702
rect 370 4600 404 4634
rect 370 4532 404 4566
rect 370 4464 404 4498
rect 370 4396 404 4430
rect 370 4328 404 4362
rect 370 4260 404 4294
rect 370 4192 404 4226
rect 370 4124 404 4158
rect 370 4056 404 4090
rect 370 3988 404 4022
rect 370 3920 404 3954
rect 370 3852 404 3886
rect 370 3784 404 3818
rect 546 4668 580 4702
rect 546 4600 580 4634
rect 546 4532 580 4566
rect 546 4464 580 4498
rect 546 4396 580 4430
rect 546 4328 580 4362
rect 546 4260 580 4294
rect 546 4192 580 4226
rect 546 4124 580 4158
rect 546 4056 580 4090
rect 546 3988 580 4022
rect 546 3920 580 3954
rect 546 3852 580 3886
rect 546 3784 580 3818
rect 370 3547 404 3581
rect 370 3479 404 3513
rect 370 3411 404 3445
rect 370 3343 404 3377
rect 370 3275 404 3309
rect 370 3207 404 3241
rect 370 3139 404 3173
rect 370 3071 404 3105
rect 370 3003 404 3037
rect 370 2935 404 2969
rect 370 2867 404 2901
rect 370 2799 404 2833
rect 370 2731 404 2765
rect 370 2663 404 2697
rect 546 3547 580 3581
rect 546 3479 580 3513
rect 546 3411 580 3445
rect 546 3343 580 3377
rect 546 3275 580 3309
rect 546 3207 580 3241
rect 546 3139 580 3173
rect 546 3071 580 3105
rect 546 3003 580 3037
rect 546 2935 580 2969
rect 546 2867 580 2901
rect 546 2799 580 2833
rect 546 2731 580 2765
rect 546 2663 580 2697
rect 370 2426 404 2460
rect 370 2358 404 2392
rect 370 2290 404 2324
rect 370 2222 404 2256
rect 370 2154 404 2188
rect 370 2086 404 2120
rect 370 2018 404 2052
rect 370 1950 404 1984
rect 370 1882 404 1916
rect 370 1814 404 1848
rect 370 1746 404 1780
rect 370 1678 404 1712
rect 370 1610 404 1644
rect 370 1542 404 1576
rect 546 2426 580 2460
rect 546 2358 580 2392
rect 546 2290 580 2324
rect 546 2222 580 2256
rect 546 2154 580 2188
rect 546 2086 580 2120
rect 546 2018 580 2052
rect 546 1950 580 1984
rect 546 1882 580 1916
rect 546 1814 580 1848
rect 546 1746 580 1780
rect 546 1678 580 1712
rect 546 1610 580 1644
rect 546 1542 580 1576
rect 370 1258 404 1292
rect 370 1190 404 1224
rect 370 1122 404 1156
rect 370 1054 404 1088
rect 370 986 404 1020
rect 370 918 404 952
rect 370 850 404 884
rect 370 782 404 816
rect 370 714 404 748
rect 370 646 404 680
rect 370 578 404 612
rect 370 510 404 544
rect 370 442 404 476
rect 370 374 404 408
rect 546 1258 580 1292
rect 546 1190 580 1224
rect 546 1122 580 1156
rect 546 1054 580 1088
rect 546 986 580 1020
rect 546 918 580 952
rect 546 850 580 884
rect 546 782 580 816
rect 546 714 580 748
rect 546 646 580 680
rect 546 578 580 612
rect 546 510 580 544
rect 546 442 580 476
rect 546 374 580 408
<< mvpsubdiff >>
rect 254 4788 278 4822
rect 312 4788 391 4822
rect 425 4788 525 4822
rect 559 4798 696 4822
rect 559 4788 662 4798
rect 254 4728 288 4788
rect 662 4729 696 4764
rect 254 4659 288 4694
rect 254 4590 288 4625
rect 254 4521 288 4556
rect 254 4452 288 4487
rect 254 4383 288 4418
rect 254 4314 288 4349
rect 254 4245 288 4280
rect 254 4176 288 4211
rect 254 4107 288 4142
rect 254 4038 288 4073
rect 254 3969 288 4004
rect 254 3900 288 3935
rect 254 3831 288 3866
rect 254 3762 288 3797
rect 254 3693 288 3728
rect 662 4660 696 4695
rect 662 4591 696 4626
rect 662 4522 696 4557
rect 662 4453 696 4488
rect 662 4384 696 4419
rect 662 4315 696 4350
rect 662 4246 696 4281
rect 662 4177 696 4212
rect 662 4108 696 4143
rect 662 4039 696 4074
rect 662 3970 696 4005
rect 662 3901 696 3936
rect 662 3832 696 3867
rect 662 3763 696 3798
rect 254 3624 288 3659
rect 662 3694 696 3729
rect 662 3625 696 3660
rect 254 3555 288 3590
rect 254 3486 288 3521
rect 254 3417 288 3452
rect 254 3348 288 3383
rect 254 3279 288 3314
rect 254 3210 288 3245
rect 254 3141 288 3176
rect 254 3072 288 3107
rect 254 3003 288 3038
rect 254 2934 288 2969
rect 254 2865 288 2900
rect 254 2796 288 2831
rect 254 2727 288 2762
rect 254 2658 288 2693
rect 254 2589 288 2624
rect 662 3556 696 3591
rect 662 3487 696 3522
rect 662 3418 696 3453
rect 662 3349 696 3384
rect 662 3280 696 3315
rect 662 3211 696 3246
rect 662 3142 696 3177
rect 662 3073 696 3108
rect 662 3004 696 3039
rect 662 2935 696 2970
rect 662 2866 696 2901
rect 662 2797 696 2832
rect 662 2728 696 2763
rect 662 2659 696 2694
rect 254 2520 288 2555
rect 254 2451 288 2486
rect 662 2590 696 2625
rect 662 2521 696 2556
rect 254 2382 288 2417
rect 254 2313 288 2348
rect 254 2244 288 2279
rect 254 2175 288 2210
rect 254 2106 288 2141
rect 254 2037 288 2072
rect 254 1968 288 2003
rect 254 1899 288 1934
rect 254 1830 288 1865
rect 254 1761 288 1796
rect 254 1692 288 1727
rect 254 1623 288 1658
rect 254 1554 288 1589
rect 254 1485 288 1520
rect 662 2452 696 2487
rect 662 2383 696 2418
rect 662 2314 696 2349
rect 662 2245 696 2280
rect 662 2176 696 2211
rect 662 2107 696 2142
rect 662 2038 696 2073
rect 662 1969 696 2004
rect 662 1900 696 1935
rect 662 1831 696 1866
rect 662 1762 696 1797
rect 662 1693 696 1728
rect 662 1624 696 1659
rect 662 1555 696 1590
rect 662 1486 696 1521
rect 254 1416 288 1451
rect 254 1347 288 1382
rect 662 1417 696 1452
rect 254 1278 288 1313
rect 254 1209 288 1244
rect 254 1140 288 1175
rect 254 1071 288 1106
rect 254 1002 288 1037
rect 254 933 288 968
rect 254 864 288 899
rect 254 795 288 830
rect 254 726 288 761
rect 254 657 288 692
rect 254 588 288 623
rect 254 519 288 554
rect 254 450 288 485
rect 254 381 288 416
rect 662 1348 696 1383
rect 662 1279 696 1314
rect 662 1210 696 1245
rect 662 1141 696 1176
rect 662 1072 696 1107
rect 662 1003 696 1038
rect 662 934 696 969
rect 662 865 696 900
rect 662 796 696 831
rect 662 727 696 762
rect 662 658 696 693
rect 662 589 696 624
rect 662 520 696 555
rect 662 451 696 486
rect 662 382 696 417
rect 254 312 288 347
rect 662 288 696 348
rect 288 278 352 288
rect 254 254 352 278
rect 386 254 423 288
rect 457 254 494 288
rect 528 254 566 288
rect 600 254 638 288
rect 672 254 696 288
<< mvnsubdiff >>
rect -852 14682 898 14686
rect -852 14648 -828 14682
rect -794 14648 -759 14682
rect -725 14648 -690 14682
rect -656 14648 -621 14682
rect -587 14648 -552 14682
rect -518 14648 -483 14682
rect -449 14648 -414 14682
rect -380 14648 -345 14682
rect -311 14648 -276 14682
rect -242 14648 -207 14682
rect -173 14648 -138 14682
rect -104 14648 -69 14682
rect -35 14648 0 14682
rect 34 14648 69 14682
rect 103 14648 138 14682
rect 172 14648 207 14682
rect 241 14648 276 14682
rect 310 14648 345 14682
rect 379 14648 414 14682
rect 448 14648 483 14682
rect 517 14648 552 14682
rect 586 14648 621 14682
rect 655 14648 690 14682
rect 724 14648 759 14682
rect 793 14648 828 14682
rect 862 14648 898 14682
rect -852 14610 898 14648
rect -852 14576 -828 14610
rect -794 14576 -759 14610
rect -725 14576 -690 14610
rect -656 14576 -621 14610
rect -587 14576 -552 14610
rect -518 14576 -483 14610
rect -449 14576 -414 14610
rect -380 14576 -345 14610
rect -311 14576 -276 14610
rect -242 14576 -207 14610
rect -173 14576 -138 14610
rect -104 14576 -69 14610
rect -35 14576 0 14610
rect 34 14576 69 14610
rect 103 14576 138 14610
rect 172 14576 207 14610
rect 241 14576 276 14610
rect 310 14576 345 14610
rect 379 14576 414 14610
rect 448 14576 483 14610
rect 517 14576 552 14610
rect 586 14576 621 14610
rect 655 14576 690 14610
rect 724 14576 759 14610
rect 793 14576 828 14610
rect 862 14576 898 14610
rect -852 14538 898 14576
rect -852 14504 -828 14538
rect -794 14504 -759 14538
rect -725 14504 -690 14538
rect -656 14504 -621 14538
rect -587 14504 -552 14538
rect -518 14504 -483 14538
rect -449 14504 -414 14538
rect -380 14504 -345 14538
rect -311 14504 -276 14538
rect -242 14504 -207 14538
rect -173 14504 -138 14538
rect -104 14504 -69 14538
rect -35 14504 0 14538
rect 34 14504 69 14538
rect 103 14504 138 14538
rect 172 14504 207 14538
rect 241 14504 276 14538
rect 310 14504 345 14538
rect 379 14504 414 14538
rect 448 14504 483 14538
rect 517 14504 552 14538
rect 586 14504 621 14538
rect 655 14504 690 14538
rect 724 14504 759 14538
rect 793 14504 828 14538
rect 862 14504 898 14538
rect -852 14466 898 14504
rect -852 14432 -828 14466
rect -794 14432 -759 14466
rect -725 14432 -690 14466
rect -656 14432 -621 14466
rect -587 14432 -552 14466
rect -518 14432 -483 14466
rect -449 14432 -414 14466
rect -380 14432 -345 14466
rect -311 14432 -276 14466
rect -242 14432 -207 14466
rect -173 14432 -138 14466
rect -104 14432 -69 14466
rect -35 14432 0 14466
rect 34 14432 69 14466
rect 103 14432 138 14466
rect 172 14432 207 14466
rect 241 14432 276 14466
rect 310 14432 345 14466
rect 379 14432 414 14466
rect 448 14432 483 14466
rect 517 14432 552 14466
rect 586 14432 621 14466
rect 655 14432 690 14466
rect 724 14432 759 14466
rect 793 14432 828 14466
rect 862 14432 898 14466
rect -852 14394 898 14432
rect -852 14360 -828 14394
rect -794 14360 -759 14394
rect -725 14360 -690 14394
rect -656 14360 -621 14394
rect -587 14360 -552 14394
rect -518 14360 -483 14394
rect -449 14360 -414 14394
rect -380 14360 -345 14394
rect -311 14360 -276 14394
rect -242 14360 -207 14394
rect -173 14360 -138 14394
rect -104 14360 -69 14394
rect -35 14360 0 14394
rect 34 14360 69 14394
rect 103 14360 138 14394
rect 172 14360 207 14394
rect 241 14360 276 14394
rect 310 14360 345 14394
rect 379 14360 414 14394
rect 448 14360 483 14394
rect 517 14360 552 14394
rect 586 14360 621 14394
rect 655 14360 690 14394
rect 724 14360 759 14394
rect 793 14360 828 14394
rect 862 14360 898 14394
rect -852 14322 898 14360
rect -852 14288 -828 14322
rect -794 14288 -759 14322
rect -725 14288 -690 14322
rect -656 14288 -621 14322
rect -587 14288 -552 14322
rect -518 14288 -483 14322
rect -449 14288 -414 14322
rect -380 14288 -345 14322
rect -311 14288 -276 14322
rect -242 14288 -207 14322
rect -173 14288 -138 14322
rect -104 14288 -69 14322
rect -35 14288 0 14322
rect 34 14288 69 14322
rect 103 14288 138 14322
rect 172 14288 207 14322
rect 241 14288 276 14322
rect 310 14288 345 14322
rect 379 14288 414 14322
rect 448 14288 483 14322
rect 517 14288 552 14322
rect 586 14288 621 14322
rect 655 14288 690 14322
rect 724 14288 759 14322
rect 793 14288 828 14322
rect 862 14288 898 14322
rect -852 14250 898 14288
rect -852 14216 -828 14250
rect -794 14216 -759 14250
rect -725 14216 -690 14250
rect -656 14216 -621 14250
rect -587 14216 -552 14250
rect -518 14216 -483 14250
rect -449 14216 -414 14250
rect -380 14216 -345 14250
rect -311 14216 -276 14250
rect -242 14216 -207 14250
rect -173 14216 -138 14250
rect -104 14216 -69 14250
rect -35 14216 0 14250
rect 34 14216 69 14250
rect 103 14216 138 14250
rect 172 14216 207 14250
rect 241 14216 276 14250
rect 310 14216 345 14250
rect 379 14216 414 14250
rect 448 14216 483 14250
rect 517 14216 552 14250
rect 586 14216 621 14250
rect 655 14216 690 14250
rect 724 14216 759 14250
rect 793 14216 828 14250
rect 862 14216 898 14250
rect -852 14178 898 14216
rect -852 14144 -828 14178
rect -794 14144 -759 14178
rect -725 14144 -690 14178
rect -656 14144 -621 14178
rect -587 14144 -552 14178
rect -518 14144 -483 14178
rect -449 14144 -414 14178
rect -380 14144 -345 14178
rect -311 14144 -276 14178
rect -242 14144 -207 14178
rect -173 14144 -138 14178
rect -104 14144 -69 14178
rect -35 14144 0 14178
rect 34 14144 69 14178
rect 103 14144 138 14178
rect 172 14144 207 14178
rect 241 14144 276 14178
rect 310 14144 345 14178
rect 379 14144 414 14178
rect 448 14144 483 14178
rect 517 14144 552 14178
rect 586 14144 621 14178
rect 655 14144 690 14178
rect 724 14144 759 14178
rect 793 14144 828 14178
rect 862 14144 898 14178
rect -852 14106 898 14144
rect -852 14072 -828 14106
rect -794 14072 -759 14106
rect -725 14072 -690 14106
rect -656 14072 -621 14106
rect -587 14072 -552 14106
rect -518 14072 -483 14106
rect -449 14072 -414 14106
rect -380 14072 -345 14106
rect -311 14072 -276 14106
rect -242 14072 -207 14106
rect -173 14072 -138 14106
rect -104 14072 -69 14106
rect -35 14072 0 14106
rect 34 14072 69 14106
rect 103 14072 138 14106
rect 172 14072 207 14106
rect 241 14072 276 14106
rect 310 14072 345 14106
rect 379 14072 414 14106
rect 448 14072 483 14106
rect 517 14072 552 14106
rect 586 14072 621 14106
rect 655 14072 690 14106
rect 724 14072 759 14106
rect 793 14072 828 14106
rect 862 14072 898 14106
rect -852 14034 898 14072
rect -852 14000 -828 14034
rect -794 14000 -759 14034
rect -725 14000 -690 14034
rect -656 14000 -621 14034
rect -587 14000 -552 14034
rect -518 14000 -483 14034
rect -449 14000 -414 14034
rect -380 14000 -345 14034
rect -311 14000 -276 14034
rect -242 14000 -207 14034
rect -173 14000 -138 14034
rect -104 14000 -69 14034
rect -35 14000 0 14034
rect 34 14000 69 14034
rect 103 14000 138 14034
rect 172 14000 207 14034
rect 241 14000 276 14034
rect 310 14000 345 14034
rect 379 14000 414 14034
rect 448 14000 483 14034
rect 517 14000 552 14034
rect 586 14000 621 14034
rect 655 14000 690 14034
rect 724 14000 759 14034
rect 793 14000 828 14034
rect 862 14000 898 14034
rect -852 13996 898 14000
rect -852 13966 20 13996
rect -852 13932 -818 13966
rect -784 13932 -748 13966
rect -714 13932 -678 13966
rect -644 13932 -608 13966
rect -574 13932 -538 13966
rect -504 13932 -468 13966
rect -434 13932 -398 13966
rect -364 13932 -328 13966
rect -294 13932 -258 13966
rect -224 13932 -188 13966
rect -154 13932 -118 13966
rect -84 13932 -48 13966
rect -14 13932 20 13966
rect -852 13898 20 13932
rect -852 13864 -818 13898
rect -784 13864 -748 13898
rect -714 13864 -678 13898
rect -644 13864 -608 13898
rect -574 13864 -538 13898
rect -504 13864 -468 13898
rect -434 13864 -398 13898
rect -364 13864 -328 13898
rect -294 13864 -258 13898
rect -224 13864 -188 13898
rect -154 13864 -118 13898
rect -84 13864 -48 13898
rect -14 13864 20 13898
rect -852 13830 20 13864
rect -852 13796 -818 13830
rect -784 13796 -748 13830
rect -714 13796 -678 13830
rect -644 13796 -608 13830
rect -574 13796 -538 13830
rect -504 13796 -468 13830
rect -434 13796 -398 13830
rect -364 13796 -328 13830
rect -294 13796 -258 13830
rect -224 13796 -188 13830
rect -154 13796 -118 13830
rect -84 13796 -48 13830
rect -14 13796 20 13830
rect -852 13762 20 13796
rect -852 13728 -818 13762
rect -784 13728 -748 13762
rect -714 13728 -678 13762
rect -644 13728 -608 13762
rect -574 13728 -538 13762
rect -504 13728 -468 13762
rect -434 13728 -398 13762
rect -364 13728 -328 13762
rect -294 13728 -258 13762
rect -224 13728 -188 13762
rect -154 13728 -118 13762
rect -84 13728 -48 13762
rect -14 13728 20 13762
rect -852 13694 20 13728
rect -852 13660 -818 13694
rect -784 13660 -748 13694
rect -714 13660 -678 13694
rect -644 13660 -608 13694
rect -574 13660 -538 13694
rect -504 13660 -468 13694
rect -434 13660 -398 13694
rect -364 13660 -328 13694
rect -294 13660 -258 13694
rect -224 13660 -188 13694
rect -154 13660 -118 13694
rect -84 13660 -48 13694
rect -14 13660 20 13694
rect -852 13626 20 13660
rect -852 13592 -818 13626
rect -784 13592 -748 13626
rect -714 13592 -678 13626
rect -644 13592 -608 13626
rect -574 13592 -538 13626
rect -504 13592 -468 13626
rect -434 13592 -398 13626
rect -364 13592 -328 13626
rect -294 13592 -258 13626
rect -224 13592 -188 13626
rect -154 13592 -118 13626
rect -84 13592 -48 13626
rect -14 13592 20 13626
rect -852 13558 20 13592
rect -852 13524 -818 13558
rect -784 13524 -748 13558
rect -714 13524 -678 13558
rect -644 13524 -608 13558
rect -574 13524 -538 13558
rect -504 13524 -468 13558
rect -434 13524 -398 13558
rect -364 13524 -328 13558
rect -294 13524 -258 13558
rect -224 13524 -188 13558
rect -154 13524 -118 13558
rect -84 13524 -48 13558
rect -14 13524 20 13558
rect -852 13490 20 13524
rect -852 13456 -818 13490
rect -784 13456 -748 13490
rect -714 13456 -678 13490
rect -644 13456 -608 13490
rect -574 13456 -538 13490
rect -504 13456 -468 13490
rect -434 13456 -398 13490
rect -364 13456 -328 13490
rect -294 13456 -258 13490
rect -224 13456 -188 13490
rect -154 13456 -118 13490
rect -84 13456 -48 13490
rect -14 13456 20 13490
rect -852 13422 20 13456
rect -852 13388 -818 13422
rect -784 13388 -748 13422
rect -714 13388 -678 13422
rect -644 13388 -608 13422
rect -574 13388 -538 13422
rect -504 13388 -468 13422
rect -434 13388 -398 13422
rect -364 13388 -328 13422
rect -294 13388 -258 13422
rect -224 13388 -188 13422
rect -154 13388 -118 13422
rect -84 13388 -48 13422
rect -14 13388 20 13422
rect -852 13354 20 13388
rect -852 13320 -818 13354
rect -784 13320 -748 13354
rect -714 13320 -678 13354
rect -644 13320 -608 13354
rect -574 13320 -538 13354
rect -504 13320 -468 13354
rect -434 13320 -398 13354
rect -364 13320 -328 13354
rect -294 13320 -258 13354
rect -224 13320 -188 13354
rect -154 13320 -118 13354
rect -84 13320 -48 13354
rect -14 13320 20 13354
rect -852 13286 20 13320
rect -852 13252 -818 13286
rect -784 13252 -748 13286
rect -714 13252 -678 13286
rect -644 13252 -608 13286
rect -574 13252 -538 13286
rect -504 13252 -468 13286
rect -434 13252 -398 13286
rect -364 13252 -328 13286
rect -294 13252 -258 13286
rect -224 13252 -188 13286
rect -154 13252 -118 13286
rect -84 13252 -48 13286
rect -14 13252 20 13286
rect -852 13218 20 13252
rect -852 13184 -818 13218
rect -784 13184 -748 13218
rect -714 13184 -678 13218
rect -644 13184 -608 13218
rect -574 13184 -538 13218
rect -504 13184 -468 13218
rect -434 13184 -398 13218
rect -364 13184 -328 13218
rect -294 13184 -258 13218
rect -224 13184 -188 13218
rect -154 13184 -118 13218
rect -84 13184 -48 13218
rect -14 13184 20 13218
rect -852 13150 20 13184
rect -852 13116 -818 13150
rect -784 13116 -748 13150
rect -714 13116 -678 13150
rect -644 13116 -608 13150
rect -574 13116 -538 13150
rect -504 13116 -468 13150
rect -434 13116 -398 13150
rect -364 13116 -328 13150
rect -294 13116 -258 13150
rect -224 13116 -188 13150
rect -154 13116 -118 13150
rect -84 13116 -48 13150
rect -14 13116 20 13150
rect -852 13082 20 13116
rect -852 13048 -818 13082
rect -784 13048 -748 13082
rect -714 13048 -678 13082
rect -644 13048 -608 13082
rect -574 13048 -538 13082
rect -504 13048 -468 13082
rect -434 13048 -398 13082
rect -364 13048 -328 13082
rect -294 13048 -258 13082
rect -224 13048 -188 13082
rect -154 13048 -118 13082
rect -84 13048 -48 13082
rect -14 13048 20 13082
rect -852 13014 20 13048
rect -852 12980 -818 13014
rect -784 12980 -748 13014
rect -714 12980 -678 13014
rect -644 12980 -608 13014
rect -574 12980 -538 13014
rect -504 12980 -468 13014
rect -434 12980 -398 13014
rect -364 12980 -328 13014
rect -294 12980 -258 13014
rect -224 12980 -188 13014
rect -154 12980 -118 13014
rect -84 12980 -48 13014
rect -14 12980 20 13014
rect -852 12946 20 12980
rect -852 12912 -818 12946
rect -784 12912 -748 12946
rect -714 12912 -678 12946
rect -644 12912 -608 12946
rect -574 12912 -538 12946
rect -504 12912 -468 12946
rect -434 12912 -398 12946
rect -364 12912 -328 12946
rect -294 12912 -258 12946
rect -224 12912 -188 12946
rect -154 12912 -118 12946
rect -84 12912 -48 12946
rect -14 12912 20 12946
rect -852 12878 20 12912
rect -852 12844 -818 12878
rect -784 12844 -748 12878
rect -714 12844 -678 12878
rect -644 12844 -608 12878
rect -574 12844 -538 12878
rect -504 12844 -468 12878
rect -434 12844 -398 12878
rect -364 12844 -328 12878
rect -294 12844 -258 12878
rect -224 12844 -188 12878
rect -154 12844 -118 12878
rect -84 12844 -48 12878
rect -14 12844 20 12878
rect -852 12810 20 12844
rect -852 12776 -818 12810
rect -784 12776 -748 12810
rect -714 12776 -678 12810
rect -644 12776 -608 12810
rect -574 12776 -538 12810
rect -504 12776 -468 12810
rect -434 12776 -398 12810
rect -364 12776 -328 12810
rect -294 12776 -258 12810
rect -224 12776 -188 12810
rect -154 12776 -118 12810
rect -84 12776 -48 12810
rect -14 12776 20 12810
rect -852 12742 20 12776
rect -852 12708 -818 12742
rect -784 12708 -748 12742
rect -714 12708 -678 12742
rect -644 12708 -608 12742
rect -574 12708 -538 12742
rect -504 12708 -468 12742
rect -434 12708 -398 12742
rect -364 12708 -328 12742
rect -294 12708 -258 12742
rect -224 12708 -188 12742
rect -154 12708 -118 12742
rect -84 12708 -48 12742
rect -14 12708 20 12742
rect -852 12674 20 12708
rect -852 12640 -818 12674
rect -784 12640 -748 12674
rect -714 12640 -678 12674
rect -644 12640 -608 12674
rect -574 12640 -538 12674
rect -504 12640 -468 12674
rect -434 12640 -398 12674
rect -364 12640 -328 12674
rect -294 12640 -258 12674
rect -224 12640 -188 12674
rect -154 12640 -118 12674
rect -84 12640 -48 12674
rect -14 12640 20 12674
rect -852 12606 20 12640
rect -852 12572 -818 12606
rect -784 12572 -748 12606
rect -714 12572 -678 12606
rect -644 12572 -608 12606
rect -574 12572 -538 12606
rect -504 12572 -468 12606
rect -434 12572 -398 12606
rect -364 12572 -328 12606
rect -294 12572 -258 12606
rect -224 12572 -188 12606
rect -154 12572 -118 12606
rect -84 12572 -48 12606
rect -14 12572 20 12606
rect -852 12538 20 12572
rect -852 12504 -818 12538
rect -784 12504 -748 12538
rect -714 12504 -678 12538
rect -644 12504 -608 12538
rect -574 12504 -538 12538
rect -504 12504 -468 12538
rect -434 12504 -398 12538
rect -364 12504 -328 12538
rect -294 12504 -258 12538
rect -224 12504 -188 12538
rect -154 12504 -118 12538
rect -84 12504 -48 12538
rect -14 12504 20 12538
rect -852 12470 20 12504
rect -852 12436 -818 12470
rect -784 12436 -748 12470
rect -714 12436 -678 12470
rect -644 12436 -608 12470
rect -574 12436 -538 12470
rect -504 12436 -468 12470
rect -434 12436 -398 12470
rect -364 12436 -328 12470
rect -294 12436 -258 12470
rect -224 12436 -188 12470
rect -154 12436 -118 12470
rect -84 12436 -48 12470
rect -14 12436 20 12470
rect -852 12402 20 12436
rect -852 12368 -818 12402
rect -784 12368 -748 12402
rect -714 12368 -678 12402
rect -644 12368 -608 12402
rect -574 12368 -538 12402
rect -504 12368 -468 12402
rect -434 12368 -398 12402
rect -364 12368 -328 12402
rect -294 12368 -258 12402
rect -224 12368 -188 12402
rect -154 12368 -118 12402
rect -84 12368 -48 12402
rect -14 12368 20 12402
rect -852 12334 20 12368
rect -852 12300 -818 12334
rect -784 12300 -748 12334
rect -714 12300 -678 12334
rect -644 12300 -608 12334
rect -574 12300 -538 12334
rect -504 12300 -468 12334
rect -434 12300 -398 12334
rect -364 12300 -328 12334
rect -294 12300 -258 12334
rect -224 12300 -188 12334
rect -154 12300 -118 12334
rect -84 12300 -48 12334
rect -14 12300 20 12334
rect -852 12266 20 12300
rect -852 12232 -818 12266
rect -784 12232 -748 12266
rect -714 12232 -678 12266
rect -644 12232 -608 12266
rect -574 12232 -538 12266
rect -504 12232 -468 12266
rect -434 12232 -398 12266
rect -364 12232 -328 12266
rect -294 12232 -258 12266
rect -224 12232 -188 12266
rect -154 12232 -118 12266
rect -84 12232 -48 12266
rect -14 12232 20 12266
rect -852 12198 20 12232
rect -852 12164 -818 12198
rect -784 12164 -748 12198
rect -714 12164 -678 12198
rect -644 12164 -608 12198
rect -574 12164 -538 12198
rect -504 12164 -468 12198
rect -434 12164 -398 12198
rect -364 12164 -328 12198
rect -294 12164 -258 12198
rect -224 12164 -188 12198
rect -154 12164 -118 12198
rect -84 12164 -48 12198
rect -14 12164 20 12198
rect -852 12160 20 12164
rect -852 12130 68 12160
rect -852 12096 -818 12130
rect -784 12096 -748 12130
rect -714 12096 -678 12130
rect -644 12096 -608 12130
rect -574 12096 -538 12130
rect -504 12096 -468 12130
rect -434 12096 -398 12130
rect -364 12096 -328 12130
rect -294 12096 -258 12130
rect -224 12096 -188 12130
rect -154 12096 -118 12130
rect -84 12096 -48 12130
rect -14 12096 68 12130
rect -852 12062 68 12096
rect -852 12028 -818 12062
rect -784 12028 -748 12062
rect -714 12028 -678 12062
rect -644 12028 -608 12062
rect -574 12028 -538 12062
rect -504 12028 -468 12062
rect -434 12028 -398 12062
rect -364 12028 -328 12062
rect -294 12028 -258 12062
rect -224 12028 -188 12062
rect -154 12028 -118 12062
rect -84 12028 -48 12062
rect -14 12028 68 12062
rect -852 11994 68 12028
rect -852 11960 -818 11994
rect -784 11960 -748 11994
rect -714 11960 -678 11994
rect -644 11960 -608 11994
rect -574 11960 -538 11994
rect -504 11960 -468 11994
rect -434 11960 -398 11994
rect -364 11960 -328 11994
rect -294 11960 -258 11994
rect -224 11960 -188 11994
rect -154 11960 -118 11994
rect -84 11960 -48 11994
rect -14 11960 68 11994
rect -852 11926 68 11960
rect -852 11892 -818 11926
rect -784 11892 -748 11926
rect -714 11892 -678 11926
rect -644 11892 -608 11926
rect -574 11892 -538 11926
rect -504 11892 -468 11926
rect -434 11892 -398 11926
rect -364 11892 -328 11926
rect -294 11892 -258 11926
rect -224 11892 -188 11926
rect -154 11892 -118 11926
rect -84 11892 -48 11926
rect -14 11892 68 11926
rect -852 11858 68 11892
rect -852 11824 -818 11858
rect -784 11824 -748 11858
rect -714 11824 -678 11858
rect -644 11824 -608 11858
rect -574 11824 -538 11858
rect -504 11824 -468 11858
rect -434 11824 -398 11858
rect -364 11824 -328 11858
rect -294 11824 -258 11858
rect -224 11824 -188 11858
rect -154 11824 -118 11858
rect -84 11824 -48 11858
rect -14 11824 68 11858
rect -852 11790 68 11824
rect -852 11756 -818 11790
rect -784 11756 -748 11790
rect -714 11756 -678 11790
rect -644 11756 -608 11790
rect -574 11756 -538 11790
rect -504 11756 -468 11790
rect -434 11756 -398 11790
rect -364 11756 -328 11790
rect -294 11756 -258 11790
rect -224 11756 -188 11790
rect -154 11756 -118 11790
rect -84 11756 -48 11790
rect -14 11756 68 11790
rect -852 11722 68 11756
rect -852 11688 -818 11722
rect -784 11688 -748 11722
rect -714 11688 -678 11722
rect -644 11688 -608 11722
rect -574 11688 -538 11722
rect -504 11688 -468 11722
rect -434 11688 -398 11722
rect -364 11688 -328 11722
rect -294 11688 -258 11722
rect -224 11688 -188 11722
rect -154 11688 -118 11722
rect -84 11688 -48 11722
rect -14 11688 68 11722
rect -852 11654 68 11688
rect -852 11620 -818 11654
rect -784 11620 -748 11654
rect -714 11620 -678 11654
rect -644 11620 -608 11654
rect -574 11620 -538 11654
rect -504 11620 -468 11654
rect -434 11620 -398 11654
rect -364 11620 -328 11654
rect -294 11620 -258 11654
rect -224 11620 -188 11654
rect -154 11620 -118 11654
rect -84 11620 -48 11654
rect -14 11620 68 11654
rect -852 11586 68 11620
rect -852 11552 -818 11586
rect -784 11552 -748 11586
rect -714 11552 -678 11586
rect -644 11552 -608 11586
rect -574 11552 -538 11586
rect -504 11552 -468 11586
rect -434 11552 -398 11586
rect -364 11552 -328 11586
rect -294 11552 -258 11586
rect -224 11552 -188 11586
rect -154 11552 -118 11586
rect -84 11552 -48 11586
rect -14 11552 68 11586
rect -852 11518 68 11552
rect -852 11484 -818 11518
rect -784 11484 -748 11518
rect -714 11484 -678 11518
rect -644 11484 -608 11518
rect -574 11484 -538 11518
rect -504 11484 -468 11518
rect -434 11484 -398 11518
rect -364 11484 -328 11518
rect -294 11484 -258 11518
rect -224 11484 -188 11518
rect -154 11484 -118 11518
rect -84 11484 -48 11518
rect -14 11484 68 11518
rect -852 11450 68 11484
rect -852 11416 -818 11450
rect -784 11416 -748 11450
rect -714 11416 -678 11450
rect -644 11416 -608 11450
rect -574 11416 -538 11450
rect -504 11416 -468 11450
rect -434 11416 -398 11450
rect -364 11416 -328 11450
rect -294 11416 -258 11450
rect -224 11416 -188 11450
rect -154 11416 -118 11450
rect -84 11416 -48 11450
rect -14 11416 68 11450
rect -852 11382 68 11416
rect -852 11348 -818 11382
rect -784 11348 -748 11382
rect -714 11348 -678 11382
rect -644 11348 -608 11382
rect -574 11348 -538 11382
rect -504 11348 -468 11382
rect -434 11348 -398 11382
rect -364 11348 -328 11382
rect -294 11348 -258 11382
rect -224 11348 -188 11382
rect -154 11348 -118 11382
rect -84 11348 -48 11382
rect -14 11348 68 11382
rect -852 11314 68 11348
rect -852 11280 -818 11314
rect -784 11280 -748 11314
rect -714 11280 -678 11314
rect -644 11280 -608 11314
rect -574 11280 -538 11314
rect -504 11280 -468 11314
rect -434 11280 -398 11314
rect -364 11280 -328 11314
rect -294 11280 -258 11314
rect -224 11280 -188 11314
rect -154 11280 -118 11314
rect -84 11280 -48 11314
rect -14 11280 68 11314
rect -852 11246 68 11280
rect -852 11212 -818 11246
rect -784 11212 -748 11246
rect -714 11212 -678 11246
rect -644 11212 -608 11246
rect -574 11212 -538 11246
rect -504 11212 -468 11246
rect -434 11212 -398 11246
rect -364 11212 -328 11246
rect -294 11212 -258 11246
rect -224 11212 -188 11246
rect -154 11212 -118 11246
rect -84 11212 -48 11246
rect -14 11212 68 11246
rect -852 11178 68 11212
rect -852 11144 -818 11178
rect -784 11144 -748 11178
rect -714 11144 -678 11178
rect -644 11144 -608 11178
rect -574 11144 -538 11178
rect -504 11144 -468 11178
rect -434 11144 -398 11178
rect -364 11144 -328 11178
rect -294 11144 -258 11178
rect -224 11144 -188 11178
rect -154 11144 -118 11178
rect -84 11144 -48 11178
rect -14 11144 68 11178
rect -852 11110 68 11144
rect -852 11076 -818 11110
rect -784 11076 -748 11110
rect -714 11076 -678 11110
rect -644 11076 -608 11110
rect -574 11076 -538 11110
rect -504 11076 -468 11110
rect -434 11076 -398 11110
rect -364 11076 -328 11110
rect -294 11076 -258 11110
rect -224 11076 -188 11110
rect -154 11076 -118 11110
rect -84 11076 -48 11110
rect -14 11076 68 11110
rect -852 11042 68 11076
rect -852 11008 -818 11042
rect -784 11008 -748 11042
rect -714 11008 -678 11042
rect -644 11008 -608 11042
rect -574 11008 -538 11042
rect -504 11008 -468 11042
rect -434 11008 -398 11042
rect -364 11008 -328 11042
rect -294 11008 -258 11042
rect -224 11008 -188 11042
rect -154 11008 -118 11042
rect -84 11008 -48 11042
rect -14 11008 68 11042
rect -852 10974 68 11008
rect -852 10940 -818 10974
rect -784 10940 -748 10974
rect -714 10940 -678 10974
rect -644 10940 -608 10974
rect -574 10940 -538 10974
rect -504 10940 -468 10974
rect -434 10940 -398 10974
rect -364 10940 -328 10974
rect -294 10940 -258 10974
rect -224 10940 -188 10974
rect -154 10940 -118 10974
rect -84 10940 -48 10974
rect -14 10940 68 10974
rect -852 10906 68 10940
rect -852 10872 -818 10906
rect -784 10872 -748 10906
rect -714 10872 -678 10906
rect -644 10872 -608 10906
rect -574 10872 -538 10906
rect -504 10872 -468 10906
rect -434 10872 -398 10906
rect -364 10872 -328 10906
rect -294 10872 -258 10906
rect -224 10872 -188 10906
rect -154 10872 -118 10906
rect -84 10872 -48 10906
rect -14 10872 68 10906
rect -852 10838 68 10872
rect -852 10804 -818 10838
rect -784 10804 -748 10838
rect -714 10804 -678 10838
rect -644 10804 -608 10838
rect -574 10804 -538 10838
rect -504 10804 -468 10838
rect -434 10804 -398 10838
rect -364 10804 -328 10838
rect -294 10804 -258 10838
rect -224 10804 -188 10838
rect -154 10804 -118 10838
rect -84 10804 -48 10838
rect -14 10804 68 10838
rect -852 10770 68 10804
rect -852 10736 -818 10770
rect -784 10736 -748 10770
rect -714 10736 -678 10770
rect -644 10736 -608 10770
rect -574 10736 -538 10770
rect -504 10736 -468 10770
rect -434 10736 -398 10770
rect -364 10736 -328 10770
rect -294 10736 -258 10770
rect -224 10736 -188 10770
rect -154 10736 -118 10770
rect -84 10736 -48 10770
rect -14 10736 68 10770
rect -852 10702 68 10736
rect -852 10668 -818 10702
rect -784 10668 -748 10702
rect -714 10668 -678 10702
rect -644 10668 -608 10702
rect -574 10668 -538 10702
rect -504 10668 -468 10702
rect -434 10668 -398 10702
rect -364 10668 -328 10702
rect -294 10668 -258 10702
rect -224 10668 -188 10702
rect -154 10668 -118 10702
rect -84 10668 -48 10702
rect -14 10668 68 10702
rect -852 10634 68 10668
rect -852 10600 -818 10634
rect -784 10600 -748 10634
rect -714 10600 -678 10634
rect -644 10600 -608 10634
rect -574 10600 -538 10634
rect -504 10600 -468 10634
rect -434 10600 -398 10634
rect -364 10600 -328 10634
rect -294 10600 -258 10634
rect -224 10600 -188 10634
rect -154 10600 -118 10634
rect -84 10600 -48 10634
rect -14 10600 68 10634
rect -852 10566 68 10600
rect -852 10532 -818 10566
rect -784 10532 -748 10566
rect -714 10532 -678 10566
rect -644 10532 -608 10566
rect -574 10532 -538 10566
rect -504 10532 -468 10566
rect -434 10532 -398 10566
rect -364 10532 -328 10566
rect -294 10532 -258 10566
rect -224 10532 -188 10566
rect -154 10532 -118 10566
rect -84 10532 -48 10566
rect -14 10532 68 10566
rect -852 10498 68 10532
rect -852 10464 -818 10498
rect -784 10464 -748 10498
rect -714 10464 -678 10498
rect -644 10464 -608 10498
rect -574 10464 -538 10498
rect -504 10464 -468 10498
rect -434 10464 -398 10498
rect -364 10464 -328 10498
rect -294 10464 -258 10498
rect -224 10464 -188 10498
rect -154 10464 -118 10498
rect -84 10464 -48 10498
rect -14 10464 68 10498
rect -852 10430 68 10464
rect -852 10396 -818 10430
rect -784 10396 -748 10430
rect -714 10396 -678 10430
rect -644 10396 -608 10430
rect -574 10396 -538 10430
rect -504 10396 -468 10430
rect -434 10396 -398 10430
rect -364 10396 -328 10430
rect -294 10396 -258 10430
rect -224 10396 -188 10430
rect -154 10396 -118 10430
rect -84 10396 -48 10430
rect -14 10396 68 10430
rect -852 10362 68 10396
rect -852 10328 -818 10362
rect -784 10328 -748 10362
rect -714 10328 -678 10362
rect -644 10328 -608 10362
rect -574 10328 -538 10362
rect -504 10328 -468 10362
rect -434 10328 -398 10362
rect -364 10328 -328 10362
rect -294 10328 -258 10362
rect -224 10328 -188 10362
rect -154 10328 -118 10362
rect -84 10328 -48 10362
rect -14 10328 68 10362
rect -852 10294 68 10328
rect -852 10260 -818 10294
rect -784 10260 -748 10294
rect -714 10260 -678 10294
rect -644 10260 -608 10294
rect -574 10260 -538 10294
rect -504 10260 -468 10294
rect -434 10260 -398 10294
rect -364 10260 -328 10294
rect -294 10260 -258 10294
rect -224 10260 -188 10294
rect -154 10260 -118 10294
rect -84 10260 -48 10294
rect -14 10260 68 10294
rect -852 10226 68 10260
rect -852 10192 -818 10226
rect -784 10192 -748 10226
rect -714 10192 -678 10226
rect -644 10192 -608 10226
rect -574 10192 -538 10226
rect -504 10192 -468 10226
rect -434 10192 -398 10226
rect -364 10192 -328 10226
rect -294 10192 -258 10226
rect -224 10192 -188 10226
rect -154 10192 -118 10226
rect -84 10192 -48 10226
rect -14 10192 68 10226
rect -852 10158 68 10192
rect -852 10124 -818 10158
rect -784 10124 -748 10158
rect -714 10124 -678 10158
rect -644 10124 -608 10158
rect -574 10124 -538 10158
rect -504 10124 -468 10158
rect -434 10124 -398 10158
rect -364 10124 -328 10158
rect -294 10124 -258 10158
rect -224 10124 -188 10158
rect -154 10124 -118 10158
rect -84 10124 -48 10158
rect -14 10124 68 10158
rect -852 10090 68 10124
rect -852 10056 -818 10090
rect -784 10056 -748 10090
rect -714 10056 -678 10090
rect -644 10056 -608 10090
rect -574 10056 -538 10090
rect -504 10056 -468 10090
rect -434 10056 -398 10090
rect -364 10056 -328 10090
rect -294 10056 -258 10090
rect -224 10056 -188 10090
rect -154 10056 -118 10090
rect -84 10056 -48 10090
rect -14 10056 68 10090
rect -852 10022 68 10056
rect -852 9988 -818 10022
rect -784 9988 -748 10022
rect -714 9988 -678 10022
rect -644 9988 -608 10022
rect -574 9988 -538 10022
rect -504 9988 -468 10022
rect -434 9988 -398 10022
rect -364 9988 -328 10022
rect -294 9988 -258 10022
rect -224 9988 -188 10022
rect -154 9988 -118 10022
rect -84 9988 -48 10022
rect -14 9988 68 10022
rect -852 9954 68 9988
rect -852 9920 -818 9954
rect -784 9920 -748 9954
rect -714 9920 -678 9954
rect -644 9920 -608 9954
rect -574 9920 -538 9954
rect -504 9920 -468 9954
rect -434 9920 -398 9954
rect -364 9920 -328 9954
rect -294 9920 -258 9954
rect -224 9920 -188 9954
rect -154 9920 -118 9954
rect -84 9920 -48 9954
rect -14 9920 68 9954
rect -852 9886 68 9920
rect -852 9852 -818 9886
rect -784 9852 -748 9886
rect -714 9852 -678 9886
rect -644 9852 -608 9886
rect -574 9852 -538 9886
rect -504 9852 -468 9886
rect -434 9852 -398 9886
rect -364 9852 -328 9886
rect -294 9852 -258 9886
rect -224 9852 -188 9886
rect -154 9852 -118 9886
rect -84 9852 -48 9886
rect -14 9852 68 9886
rect -852 9818 68 9852
rect -852 9784 -818 9818
rect -784 9784 -748 9818
rect -714 9784 -678 9818
rect -644 9784 -608 9818
rect -574 9784 -538 9818
rect -504 9784 -468 9818
rect -434 9784 -398 9818
rect -364 9784 -328 9818
rect -294 9784 -258 9818
rect -224 9784 -188 9818
rect -154 9784 -118 9818
rect -84 9784 -48 9818
rect -14 9784 68 9818
rect -852 9750 68 9784
rect -852 9716 -818 9750
rect -784 9716 -748 9750
rect -714 9716 -678 9750
rect -644 9716 -608 9750
rect -574 9716 -538 9750
rect -504 9716 -468 9750
rect -434 9716 -398 9750
rect -364 9716 -328 9750
rect -294 9716 -258 9750
rect -224 9716 -188 9750
rect -154 9716 -118 9750
rect -84 9716 -48 9750
rect -14 9716 68 9750
rect -852 9682 68 9716
rect -852 9648 -818 9682
rect -784 9648 -748 9682
rect -714 9648 -678 9682
rect -644 9648 -608 9682
rect -574 9648 -538 9682
rect -504 9648 -468 9682
rect -434 9648 -398 9682
rect -364 9648 -328 9682
rect -294 9648 -258 9682
rect -224 9648 -188 9682
rect -154 9648 -118 9682
rect -84 9648 -48 9682
rect -14 9648 68 9682
rect -852 9614 68 9648
rect -852 9580 -818 9614
rect -784 9580 -748 9614
rect -714 9580 -678 9614
rect -644 9580 -608 9614
rect -574 9580 -538 9614
rect -504 9580 -468 9614
rect -434 9580 -398 9614
rect -364 9580 -328 9614
rect -294 9580 -258 9614
rect -224 9580 -188 9614
rect -154 9580 -118 9614
rect -84 9580 -48 9614
rect -14 9580 68 9614
rect -852 9546 68 9580
rect -852 9512 -818 9546
rect -784 9512 -748 9546
rect -714 9512 -678 9546
rect -644 9512 -608 9546
rect -574 9512 -538 9546
rect -504 9512 -468 9546
rect -434 9512 -398 9546
rect -364 9512 -328 9546
rect -294 9512 -258 9546
rect -224 9512 -188 9546
rect -154 9512 -118 9546
rect -84 9512 -48 9546
rect -14 9512 68 9546
rect -852 9478 68 9512
rect -852 9444 -818 9478
rect -784 9444 -748 9478
rect -714 9444 -678 9478
rect -644 9444 -608 9478
rect -574 9444 -538 9478
rect -504 9444 -468 9478
rect -434 9444 -398 9478
rect -364 9444 -328 9478
rect -294 9444 -258 9478
rect -224 9444 -188 9478
rect -154 9444 -118 9478
rect -84 9444 -48 9478
rect -14 9444 68 9478
rect -852 9410 68 9444
rect -852 9376 -818 9410
rect -784 9376 -748 9410
rect -714 9376 -678 9410
rect -644 9376 -608 9410
rect -574 9376 -538 9410
rect -504 9376 -468 9410
rect -434 9376 -398 9410
rect -364 9376 -328 9410
rect -294 9376 -258 9410
rect -224 9376 -188 9410
rect -154 9376 -118 9410
rect -84 9376 -48 9410
rect -14 9376 68 9410
rect -852 9342 68 9376
rect -852 9308 -818 9342
rect -784 9308 -748 9342
rect -714 9308 -678 9342
rect -644 9308 -608 9342
rect -574 9308 -538 9342
rect -504 9308 -468 9342
rect -434 9308 -398 9342
rect -364 9308 -328 9342
rect -294 9308 -258 9342
rect -224 9308 -188 9342
rect -154 9308 -118 9342
rect -84 9308 -48 9342
rect -14 9308 68 9342
rect -852 9274 68 9308
rect -852 9240 -818 9274
rect -784 9240 -748 9274
rect -714 9240 -678 9274
rect -644 9240 -608 9274
rect -574 9240 -538 9274
rect -504 9240 -468 9274
rect -434 9240 -398 9274
rect -364 9240 -328 9274
rect -294 9240 -258 9274
rect -224 9240 -188 9274
rect -154 9240 -118 9274
rect -84 9240 -48 9274
rect -14 9240 68 9274
rect -852 9206 68 9240
rect -852 9172 -818 9206
rect -784 9172 -748 9206
rect -714 9172 -678 9206
rect -644 9172 -608 9206
rect -574 9172 -538 9206
rect -504 9172 -468 9206
rect -434 9172 -398 9206
rect -364 9172 -328 9206
rect -294 9172 -258 9206
rect -224 9172 -188 9206
rect -154 9172 -118 9206
rect -84 9172 -48 9206
rect -14 9172 68 9206
rect -852 9138 68 9172
rect -852 9104 -818 9138
rect -784 9104 -748 9138
rect -714 9104 -678 9138
rect -644 9104 -608 9138
rect -574 9104 -538 9138
rect -504 9104 -468 9138
rect -434 9104 -398 9138
rect -364 9104 -328 9138
rect -294 9104 -258 9138
rect -224 9104 -188 9138
rect -154 9104 -118 9138
rect -84 9104 -48 9138
rect -14 9104 68 9138
rect -852 9070 68 9104
rect -852 9036 -818 9070
rect -784 9036 -748 9070
rect -714 9036 -678 9070
rect -644 9036 -608 9070
rect -574 9036 -538 9070
rect -504 9036 -468 9070
rect -434 9036 -398 9070
rect -364 9036 -328 9070
rect -294 9036 -258 9070
rect -224 9036 -188 9070
rect -154 9036 -118 9070
rect -84 9036 -48 9070
rect -14 9036 68 9070
rect -852 9002 68 9036
rect -852 8968 -818 9002
rect -784 8968 -748 9002
rect -714 8968 -678 9002
rect -644 8968 -608 9002
rect -574 8968 -538 9002
rect -504 8968 -468 9002
rect -434 8968 -398 9002
rect -364 8968 -328 9002
rect -294 8968 -258 9002
rect -224 8968 -188 9002
rect -154 8968 -118 9002
rect -84 8968 -48 9002
rect -14 8968 68 9002
rect -852 8934 68 8968
rect -852 8900 -818 8934
rect -784 8900 -748 8934
rect -714 8900 -678 8934
rect -644 8900 -608 8934
rect -574 8900 -538 8934
rect -504 8900 -468 8934
rect -434 8900 -398 8934
rect -364 8900 -328 8934
rect -294 8900 -258 8934
rect -224 8900 -188 8934
rect -154 8900 -118 8934
rect -84 8900 -48 8934
rect -14 8900 68 8934
rect -852 8866 68 8900
rect -852 8832 -818 8866
rect -784 8832 -748 8866
rect -714 8832 -678 8866
rect -644 8832 -608 8866
rect -574 8832 -538 8866
rect -504 8832 -468 8866
rect -434 8832 -398 8866
rect -364 8832 -328 8866
rect -294 8832 -258 8866
rect -224 8832 -188 8866
rect -154 8832 -118 8866
rect -84 8832 -48 8866
rect -14 8832 68 8866
rect -852 8798 68 8832
rect -852 8764 -818 8798
rect -784 8764 -748 8798
rect -714 8764 -678 8798
rect -644 8764 -608 8798
rect -574 8764 -538 8798
rect -504 8764 -468 8798
rect -434 8764 -398 8798
rect -364 8764 -328 8798
rect -294 8764 -258 8798
rect -224 8764 -188 8798
rect -154 8764 -118 8798
rect -84 8764 -48 8798
rect -14 8764 68 8798
rect -852 8730 68 8764
rect -852 8696 -818 8730
rect -784 8696 -748 8730
rect -714 8696 -678 8730
rect -644 8696 -608 8730
rect -574 8696 -538 8730
rect -504 8696 -468 8730
rect -434 8696 -398 8730
rect -364 8696 -328 8730
rect -294 8696 -258 8730
rect -224 8696 -188 8730
rect -154 8696 -118 8730
rect -84 8696 -48 8730
rect -14 8696 68 8730
rect -852 8662 68 8696
rect -852 8628 -818 8662
rect -784 8628 -748 8662
rect -714 8628 -678 8662
rect -644 8628 -608 8662
rect -574 8628 -538 8662
rect -504 8628 -468 8662
rect -434 8628 -398 8662
rect -364 8628 -328 8662
rect -294 8628 -258 8662
rect -224 8628 -188 8662
rect -154 8628 -118 8662
rect -84 8628 -48 8662
rect -14 8628 68 8662
rect -852 8594 68 8628
rect -852 8560 -818 8594
rect -784 8560 -748 8594
rect -714 8560 -678 8594
rect -644 8560 -608 8594
rect -574 8560 -538 8594
rect -504 8560 -468 8594
rect -434 8560 -398 8594
rect -364 8560 -328 8594
rect -294 8560 -258 8594
rect -224 8560 -188 8594
rect -154 8560 -118 8594
rect -84 8560 -48 8594
rect -14 8560 68 8594
rect -852 8526 68 8560
rect -852 8492 -818 8526
rect -784 8492 -748 8526
rect -714 8492 -678 8526
rect -644 8492 -608 8526
rect -574 8492 -538 8526
rect -504 8492 -468 8526
rect -434 8492 -398 8526
rect -364 8492 -328 8526
rect -294 8492 -258 8526
rect -224 8492 -188 8526
rect -154 8492 -118 8526
rect -84 8492 -48 8526
rect -14 8492 68 8526
rect -852 8458 68 8492
rect -852 8424 -818 8458
rect -784 8424 -748 8458
rect -714 8424 -678 8458
rect -644 8424 -608 8458
rect -574 8424 -538 8458
rect -504 8424 -468 8458
rect -434 8424 -398 8458
rect -364 8424 -328 8458
rect -294 8424 -258 8458
rect -224 8424 -188 8458
rect -154 8424 -118 8458
rect -84 8424 -48 8458
rect -14 8424 68 8458
rect -852 8390 68 8424
rect -852 8356 -818 8390
rect -784 8356 -748 8390
rect -714 8356 -678 8390
rect -644 8356 -608 8390
rect -574 8356 -538 8390
rect -504 8356 -468 8390
rect -434 8356 -398 8390
rect -364 8356 -328 8390
rect -294 8356 -258 8390
rect -224 8356 -188 8390
rect -154 8356 -118 8390
rect -84 8356 -48 8390
rect -14 8356 68 8390
rect -852 8322 68 8356
rect -852 8288 -818 8322
rect -784 8288 -748 8322
rect -714 8288 -678 8322
rect -644 8288 -608 8322
rect -574 8288 -538 8322
rect -504 8288 -468 8322
rect -434 8288 -398 8322
rect -364 8288 -328 8322
rect -294 8288 -258 8322
rect -224 8288 -188 8322
rect -154 8288 -118 8322
rect -84 8288 -48 8322
rect -14 8288 68 8322
rect -852 8254 68 8288
rect -852 8220 -818 8254
rect -784 8220 -748 8254
rect -714 8220 -678 8254
rect -644 8220 -608 8254
rect -574 8220 -538 8254
rect -504 8220 -468 8254
rect -434 8220 -398 8254
rect -364 8220 -328 8254
rect -294 8220 -258 8254
rect -224 8220 -188 8254
rect -154 8220 -118 8254
rect -84 8220 -48 8254
rect -14 8220 68 8254
rect -852 8186 68 8220
rect -852 8152 -818 8186
rect -784 8152 -748 8186
rect -714 8152 -678 8186
rect -644 8152 -608 8186
rect -574 8152 -538 8186
rect -504 8152 -468 8186
rect -434 8152 -398 8186
rect -364 8152 -328 8186
rect -294 8152 -258 8186
rect -224 8152 -188 8186
rect -154 8152 -118 8186
rect -84 8152 -48 8186
rect -14 8152 68 8186
rect -852 8118 68 8152
rect -852 8084 -818 8118
rect -784 8084 -748 8118
rect -714 8084 -678 8118
rect -644 8084 -608 8118
rect -574 8084 -538 8118
rect -504 8084 -468 8118
rect -434 8084 -398 8118
rect -364 8084 -328 8118
rect -294 8084 -258 8118
rect -224 8084 -188 8118
rect -154 8084 -118 8118
rect -84 8084 -48 8118
rect -14 8084 68 8118
rect -852 8050 68 8084
rect -852 8016 -818 8050
rect -784 8016 -748 8050
rect -714 8016 -678 8050
rect -644 8016 -608 8050
rect -574 8016 -538 8050
rect -504 8016 -468 8050
rect -434 8016 -398 8050
rect -364 8016 -328 8050
rect -294 8016 -258 8050
rect -224 8016 -188 8050
rect -154 8016 -118 8050
rect -84 8016 -48 8050
rect -14 8016 68 8050
rect -852 7982 68 8016
rect -852 7948 -818 7982
rect -784 7948 -748 7982
rect -714 7948 -678 7982
rect -644 7948 -608 7982
rect -574 7948 -538 7982
rect -504 7948 -468 7982
rect -434 7948 -398 7982
rect -364 7948 -328 7982
rect -294 7948 -258 7982
rect -224 7948 -188 7982
rect -154 7948 -118 7982
rect -84 7948 -48 7982
rect -14 7948 68 7982
rect -852 7914 68 7948
rect -852 7880 -818 7914
rect -784 7880 -748 7914
rect -714 7880 -678 7914
rect -644 7880 -608 7914
rect -574 7880 -538 7914
rect -504 7880 -468 7914
rect -434 7880 -398 7914
rect -364 7880 -328 7914
rect -294 7880 -258 7914
rect -224 7880 -188 7914
rect -154 7880 -118 7914
rect -84 7880 -48 7914
rect -14 7880 68 7914
rect -852 7846 68 7880
rect -852 7812 -818 7846
rect -784 7812 -748 7846
rect -714 7812 -678 7846
rect -644 7812 -608 7846
rect -574 7812 -538 7846
rect -504 7812 -468 7846
rect -434 7812 -398 7846
rect -364 7812 -328 7846
rect -294 7812 -258 7846
rect -224 7812 -188 7846
rect -154 7812 -118 7846
rect -84 7812 -48 7846
rect -14 7812 68 7846
rect -852 7778 68 7812
rect -852 7744 -818 7778
rect -784 7744 -748 7778
rect -714 7744 -678 7778
rect -644 7744 -608 7778
rect -574 7744 -538 7778
rect -504 7744 -468 7778
rect -434 7744 -398 7778
rect -364 7744 -328 7778
rect -294 7744 -258 7778
rect -224 7744 -188 7778
rect -154 7744 -118 7778
rect -84 7744 -48 7778
rect -14 7744 68 7778
rect -852 7710 68 7744
rect -852 7676 -818 7710
rect -784 7676 -748 7710
rect -714 7676 -678 7710
rect -644 7676 -608 7710
rect -574 7676 -538 7710
rect -504 7676 -468 7710
rect -434 7676 -398 7710
rect -364 7676 -328 7710
rect -294 7676 -258 7710
rect -224 7676 -188 7710
rect -154 7676 -118 7710
rect -84 7676 -48 7710
rect -14 7676 68 7710
rect -852 7642 68 7676
rect -852 7608 -818 7642
rect -784 7608 -748 7642
rect -714 7608 -678 7642
rect -644 7608 -608 7642
rect -574 7608 -538 7642
rect -504 7608 -468 7642
rect -434 7608 -398 7642
rect -364 7608 -328 7642
rect -294 7608 -258 7642
rect -224 7608 -188 7642
rect -154 7608 -118 7642
rect -84 7608 -48 7642
rect -14 7608 68 7642
rect -852 7574 68 7608
rect -852 7540 -818 7574
rect -784 7540 -748 7574
rect -714 7540 -678 7574
rect -644 7540 -608 7574
rect -574 7540 -538 7574
rect -504 7540 -468 7574
rect -434 7540 -398 7574
rect -364 7540 -328 7574
rect -294 7540 -258 7574
rect -224 7540 -188 7574
rect -154 7540 -118 7574
rect -84 7540 -48 7574
rect -14 7540 68 7574
rect -852 7506 68 7540
rect -852 7472 -818 7506
rect -784 7472 -748 7506
rect -714 7472 -678 7506
rect -644 7472 -608 7506
rect -574 7472 -538 7506
rect -504 7472 -468 7506
rect -434 7472 -398 7506
rect -364 7472 -328 7506
rect -294 7472 -258 7506
rect -224 7472 -188 7506
rect -154 7472 -118 7506
rect -84 7472 -48 7506
rect -14 7472 68 7506
rect -852 7438 68 7472
rect -852 7404 -818 7438
rect -784 7404 -748 7438
rect -714 7404 -678 7438
rect -644 7404 -608 7438
rect -574 7404 -538 7438
rect -504 7404 -468 7438
rect -434 7404 -398 7438
rect -364 7404 -328 7438
rect -294 7404 -258 7438
rect -224 7404 -188 7438
rect -154 7404 -118 7438
rect -84 7404 -48 7438
rect -14 7404 68 7438
rect -852 7370 68 7404
rect -852 7336 -818 7370
rect -784 7336 -748 7370
rect -714 7336 -678 7370
rect -644 7336 -608 7370
rect -574 7336 -538 7370
rect -504 7336 -468 7370
rect -434 7336 -398 7370
rect -364 7336 -328 7370
rect -294 7336 -258 7370
rect -224 7336 -188 7370
rect -154 7336 -118 7370
rect -84 7336 -48 7370
rect -14 7336 68 7370
rect -852 7302 68 7336
rect -852 7268 -818 7302
rect -784 7268 -748 7302
rect -714 7268 -678 7302
rect -644 7268 -608 7302
rect -574 7268 -538 7302
rect -504 7268 -468 7302
rect -434 7268 -398 7302
rect -364 7268 -328 7302
rect -294 7268 -258 7302
rect -224 7268 -188 7302
rect -154 7268 -118 7302
rect -84 7268 -48 7302
rect -14 7268 68 7302
rect -852 7234 68 7268
rect -852 7200 -818 7234
rect -784 7200 -748 7234
rect -714 7200 -678 7234
rect -644 7200 -608 7234
rect -574 7200 -538 7234
rect -504 7200 -468 7234
rect -434 7200 -398 7234
rect -364 7200 -328 7234
rect -294 7200 -258 7234
rect -224 7200 -188 7234
rect -154 7200 -118 7234
rect -84 7200 -48 7234
rect -14 7200 68 7234
rect -852 7166 68 7200
rect -852 7132 -818 7166
rect -784 7132 -748 7166
rect -714 7132 -678 7166
rect -644 7132 -608 7166
rect -574 7132 -538 7166
rect -504 7132 -468 7166
rect -434 7132 -398 7166
rect -364 7132 -328 7166
rect -294 7132 -258 7166
rect -224 7132 -188 7166
rect -154 7132 -118 7166
rect -84 7132 -48 7166
rect -14 7132 68 7166
rect -852 7098 68 7132
rect -852 7064 -818 7098
rect -784 7064 -748 7098
rect -714 7064 -678 7098
rect -644 7064 -608 7098
rect -574 7064 -538 7098
rect -504 7064 -468 7098
rect -434 7064 -398 7098
rect -364 7064 -328 7098
rect -294 7064 -258 7098
rect -224 7064 -188 7098
rect -154 7064 -118 7098
rect -84 7064 -48 7098
rect -14 7064 68 7098
rect -852 7030 68 7064
rect -852 6996 -818 7030
rect -784 6996 -748 7030
rect -714 6996 -678 7030
rect -644 6996 -608 7030
rect -574 6996 -538 7030
rect -504 6996 -468 7030
rect -434 6996 -398 7030
rect -364 6996 -328 7030
rect -294 6996 -258 7030
rect -224 6996 -188 7030
rect -154 6996 -118 7030
rect -84 6996 -48 7030
rect -14 6996 68 7030
rect -852 6962 68 6996
rect -852 6928 -818 6962
rect -784 6928 -748 6962
rect -714 6928 -678 6962
rect -644 6928 -608 6962
rect -574 6928 -538 6962
rect -504 6928 -468 6962
rect -434 6928 -398 6962
rect -364 6928 -328 6962
rect -294 6928 -258 6962
rect -224 6928 -188 6962
rect -154 6928 -118 6962
rect -84 6928 -48 6962
rect -14 6928 68 6962
rect -852 6894 68 6928
rect -852 6860 -818 6894
rect -784 6860 -748 6894
rect -714 6860 -678 6894
rect -644 6860 -608 6894
rect -574 6860 -538 6894
rect -504 6860 -468 6894
rect -434 6860 -398 6894
rect -364 6860 -328 6894
rect -294 6860 -258 6894
rect -224 6860 -188 6894
rect -154 6860 -118 6894
rect -84 6860 -48 6894
rect -14 6860 68 6894
rect -852 6826 68 6860
rect -852 6792 -818 6826
rect -784 6792 -748 6826
rect -714 6792 -678 6826
rect -644 6792 -608 6826
rect -574 6792 -538 6826
rect -504 6792 -468 6826
rect -434 6792 -398 6826
rect -364 6792 -328 6826
rect -294 6792 -258 6826
rect -224 6792 -188 6826
rect -154 6792 -118 6826
rect -84 6792 -48 6826
rect -14 6792 68 6826
rect -852 6758 68 6792
rect -852 6724 -818 6758
rect -784 6724 -748 6758
rect -714 6724 -678 6758
rect -644 6724 -608 6758
rect -574 6724 -538 6758
rect -504 6724 -468 6758
rect -434 6724 -398 6758
rect -364 6724 -328 6758
rect -294 6724 -258 6758
rect -224 6724 -188 6758
rect -154 6724 -118 6758
rect -84 6724 -48 6758
rect -14 6724 68 6758
rect -852 6690 68 6724
rect -852 6656 -818 6690
rect -784 6656 -748 6690
rect -714 6656 -678 6690
rect -644 6656 -608 6690
rect -574 6656 -538 6690
rect -504 6656 -468 6690
rect -434 6656 -398 6690
rect -364 6656 -328 6690
rect -294 6656 -258 6690
rect -224 6656 -188 6690
rect -154 6656 -118 6690
rect -84 6656 -48 6690
rect -14 6656 68 6690
rect -852 6622 68 6656
rect -852 6588 -818 6622
rect -784 6588 -748 6622
rect -714 6588 -678 6622
rect -644 6588 -608 6622
rect -574 6588 -538 6622
rect -504 6588 -468 6622
rect -434 6588 -398 6622
rect -364 6588 -328 6622
rect -294 6588 -258 6622
rect -224 6588 -188 6622
rect -154 6588 -118 6622
rect -84 6588 -48 6622
rect -14 6588 68 6622
rect -852 6554 68 6588
rect -852 6520 -818 6554
rect -784 6520 -748 6554
rect -714 6520 -678 6554
rect -644 6520 -608 6554
rect -574 6520 -538 6554
rect -504 6520 -468 6554
rect -434 6520 -398 6554
rect -364 6520 -328 6554
rect -294 6520 -258 6554
rect -224 6520 -188 6554
rect -154 6520 -118 6554
rect -84 6520 -48 6554
rect -14 6520 68 6554
rect -852 6486 68 6520
rect -852 6452 -818 6486
rect -784 6452 -748 6486
rect -714 6452 -678 6486
rect -644 6452 -608 6486
rect -574 6452 -538 6486
rect -504 6452 -468 6486
rect -434 6452 -398 6486
rect -364 6452 -328 6486
rect -294 6452 -258 6486
rect -224 6452 -188 6486
rect -154 6452 -118 6486
rect -84 6452 -48 6486
rect -14 6452 68 6486
rect -852 6418 68 6452
rect -852 6384 -818 6418
rect -784 6384 -748 6418
rect -714 6384 -678 6418
rect -644 6384 -608 6418
rect -574 6384 -538 6418
rect -504 6384 -468 6418
rect -434 6384 -398 6418
rect -364 6384 -328 6418
rect -294 6384 -258 6418
rect -224 6384 -188 6418
rect -154 6384 -118 6418
rect -84 6384 -48 6418
rect -14 6384 68 6418
rect -852 6350 68 6384
rect -852 6316 -818 6350
rect -784 6316 -748 6350
rect -714 6316 -678 6350
rect -644 6316 -608 6350
rect -574 6316 -538 6350
rect -504 6316 -468 6350
rect -434 6316 -398 6350
rect -364 6316 -328 6350
rect -294 6316 -258 6350
rect -224 6316 -188 6350
rect -154 6316 -118 6350
rect -84 6316 -48 6350
rect -14 6316 68 6350
rect -852 6282 68 6316
rect -852 6248 -818 6282
rect -784 6248 -748 6282
rect -714 6248 -678 6282
rect -644 6248 -608 6282
rect -574 6248 -538 6282
rect -504 6248 -468 6282
rect -434 6248 -398 6282
rect -364 6248 -328 6282
rect -294 6248 -258 6282
rect -224 6248 -188 6282
rect -154 6248 -118 6282
rect -84 6248 -48 6282
rect -14 6248 68 6282
rect -852 6214 68 6248
rect -852 6180 -818 6214
rect -784 6180 -748 6214
rect -714 6180 -678 6214
rect -644 6180 -608 6214
rect -574 6180 -538 6214
rect -504 6180 -468 6214
rect -434 6180 -398 6214
rect -364 6180 -328 6214
rect -294 6180 -258 6214
rect -224 6180 -188 6214
rect -154 6180 -118 6214
rect -84 6180 -48 6214
rect -14 6180 68 6214
rect -852 6146 68 6180
rect -852 6112 -818 6146
rect -784 6112 -748 6146
rect -714 6112 -678 6146
rect -644 6112 -608 6146
rect -574 6112 -538 6146
rect -504 6112 -468 6146
rect -434 6112 -398 6146
rect -364 6112 -328 6146
rect -294 6112 -258 6146
rect -224 6112 -188 6146
rect -154 6112 -118 6146
rect -84 6112 -48 6146
rect -14 6112 68 6146
rect -852 6078 68 6112
rect -852 6044 -818 6078
rect -784 6044 -748 6078
rect -714 6044 -678 6078
rect -644 6044 -608 6078
rect -574 6044 -538 6078
rect -504 6044 -468 6078
rect -434 6044 -398 6078
rect -364 6044 -328 6078
rect -294 6044 -258 6078
rect -224 6044 -188 6078
rect -154 6044 -118 6078
rect -84 6044 -48 6078
rect -14 6044 68 6078
rect -852 6010 68 6044
rect -852 5976 -818 6010
rect -784 5976 -748 6010
rect -714 5976 -678 6010
rect -644 5976 -608 6010
rect -574 5976 -538 6010
rect -504 5976 -468 6010
rect -434 5976 -398 6010
rect -364 5976 -328 6010
rect -294 5976 -258 6010
rect -224 5976 -188 6010
rect -154 5976 -118 6010
rect -84 5976 -48 6010
rect -14 5976 68 6010
rect -852 5942 68 5976
rect -852 5908 -818 5942
rect -784 5908 -748 5942
rect -714 5908 -678 5942
rect -644 5908 -608 5942
rect -574 5908 -538 5942
rect -504 5908 -468 5942
rect -434 5908 -398 5942
rect -364 5908 -328 5942
rect -294 5908 -258 5942
rect -224 5908 -188 5942
rect -154 5908 -118 5942
rect -84 5908 -48 5942
rect -14 5908 68 5942
rect -852 5874 68 5908
rect -852 5840 -818 5874
rect -784 5840 -748 5874
rect -714 5840 -678 5874
rect -644 5840 -608 5874
rect -574 5840 -538 5874
rect -504 5840 -468 5874
rect -434 5840 -398 5874
rect -364 5840 -328 5874
rect -294 5840 -258 5874
rect -224 5840 -188 5874
rect -154 5840 -118 5874
rect -84 5840 -48 5874
rect -14 5840 68 5874
rect -852 5806 68 5840
rect -852 5772 -818 5806
rect -784 5772 -748 5806
rect -714 5772 -678 5806
rect -644 5772 -608 5806
rect -574 5772 -538 5806
rect -504 5772 -468 5806
rect -434 5772 -398 5806
rect -364 5772 -328 5806
rect -294 5772 -258 5806
rect -224 5772 -188 5806
rect -154 5772 -118 5806
rect -84 5772 -48 5806
rect -14 5772 68 5806
rect -852 5738 68 5772
rect -852 5704 -818 5738
rect -784 5704 -748 5738
rect -714 5704 -678 5738
rect -644 5704 -608 5738
rect -574 5704 -538 5738
rect -504 5704 -468 5738
rect -434 5704 -398 5738
rect -364 5704 -328 5738
rect -294 5704 -258 5738
rect -224 5704 -188 5738
rect -154 5704 -118 5738
rect -84 5704 -48 5738
rect -14 5704 68 5738
rect -852 5670 68 5704
rect -852 5636 -818 5670
rect -784 5636 -748 5670
rect -714 5636 -678 5670
rect -644 5636 -608 5670
rect -574 5636 -538 5670
rect -504 5636 -468 5670
rect -434 5636 -398 5670
rect -364 5636 -328 5670
rect -294 5636 -258 5670
rect -224 5636 -188 5670
rect -154 5636 -118 5670
rect -84 5636 -48 5670
rect -14 5636 68 5670
rect -852 5602 68 5636
rect -852 5568 -818 5602
rect -784 5568 -748 5602
rect -714 5568 -678 5602
rect -644 5568 -608 5602
rect -574 5568 -538 5602
rect -504 5568 -468 5602
rect -434 5568 -398 5602
rect -364 5568 -328 5602
rect -294 5568 -258 5602
rect -224 5568 -188 5602
rect -154 5568 -118 5602
rect -84 5568 -48 5602
rect -14 5568 68 5602
rect -852 5534 68 5568
rect -852 5500 -818 5534
rect -784 5500 -748 5534
rect -714 5500 -678 5534
rect -644 5500 -608 5534
rect -574 5500 -538 5534
rect -504 5500 -468 5534
rect -434 5500 -398 5534
rect -364 5500 -328 5534
rect -294 5500 -258 5534
rect -224 5500 -188 5534
rect -154 5500 -118 5534
rect -84 5500 -48 5534
rect -14 5500 68 5534
rect -852 5466 68 5500
rect -852 5432 -818 5466
rect -784 5432 -748 5466
rect -714 5432 -678 5466
rect -644 5432 -608 5466
rect -574 5432 -538 5466
rect -504 5432 -468 5466
rect -434 5432 -398 5466
rect -364 5432 -328 5466
rect -294 5432 -258 5466
rect -224 5432 -188 5466
rect -154 5432 -118 5466
rect -84 5432 -48 5466
rect -14 5432 68 5466
rect -852 5398 68 5432
rect -852 5364 -818 5398
rect -784 5364 -748 5398
rect -714 5364 -678 5398
rect -644 5364 -608 5398
rect -574 5364 -538 5398
rect -504 5364 -468 5398
rect -434 5364 -398 5398
rect -364 5364 -328 5398
rect -294 5364 -258 5398
rect -224 5364 -188 5398
rect -154 5364 -118 5398
rect -84 5364 -48 5398
rect -14 5364 68 5398
rect -852 5330 68 5364
rect -852 5296 -818 5330
rect -784 5296 -748 5330
rect -714 5296 -678 5330
rect -644 5296 -608 5330
rect -574 5296 -538 5330
rect -504 5296 -468 5330
rect -434 5296 -398 5330
rect -364 5296 -328 5330
rect -294 5296 -258 5330
rect -224 5296 -188 5330
rect -154 5296 -118 5330
rect -84 5296 -48 5330
rect -14 5296 68 5330
rect -852 5262 68 5296
rect -852 5228 -818 5262
rect -784 5228 -748 5262
rect -714 5228 -678 5262
rect -644 5228 -608 5262
rect -574 5228 -538 5262
rect -504 5228 -468 5262
rect -434 5228 -398 5262
rect -364 5228 -328 5262
rect -294 5228 -258 5262
rect -224 5228 -188 5262
rect -154 5228 -118 5262
rect -84 5228 -48 5262
rect -14 5228 68 5262
rect -852 5194 68 5228
rect -852 5160 -818 5194
rect -784 5160 -748 5194
rect -714 5160 -678 5194
rect -644 5160 -608 5194
rect -574 5160 -538 5194
rect -504 5160 -468 5194
rect -434 5160 -398 5194
rect -364 5160 -328 5194
rect -294 5160 -258 5194
rect -224 5160 -188 5194
rect -154 5160 -118 5194
rect -84 5160 -48 5194
rect -14 5160 68 5194
rect -852 5126 68 5160
rect -852 5092 -818 5126
rect -784 5092 -748 5126
rect -714 5092 -678 5126
rect -644 5092 -608 5126
rect -574 5092 -538 5126
rect -504 5092 -468 5126
rect -434 5092 -398 5126
rect -364 5092 -328 5126
rect -294 5092 -258 5126
rect -224 5092 -188 5126
rect -154 5092 -118 5126
rect -84 5092 -48 5126
rect -14 5092 68 5126
rect -852 5058 68 5092
rect -852 5024 -818 5058
rect -784 5024 -748 5058
rect -714 5024 -678 5058
rect -644 5024 -608 5058
rect -574 5024 -538 5058
rect -504 5024 -468 5058
rect -434 5024 -398 5058
rect -364 5024 -328 5058
rect -294 5024 -258 5058
rect -224 5024 -188 5058
rect -154 5024 -118 5058
rect -84 5024 -48 5058
rect -14 5024 68 5058
rect -852 5010 68 5024
rect -852 4990 882 5010
rect -852 4956 -818 4990
rect -784 4956 -748 4990
rect -714 4956 -678 4990
rect -644 4956 -608 4990
rect -574 4956 -538 4990
rect -504 4956 -468 4990
rect -434 4956 -398 4990
rect -364 4956 -328 4990
rect -294 4956 -258 4990
rect -224 4956 -188 4990
rect -154 4956 -118 4990
rect -84 4956 -48 4990
rect -14 4986 882 4990
rect -14 4956 68 4986
rect -852 4952 68 4956
rect 102 4976 882 4986
rect -852 4922 102 4952
rect -852 4888 -818 4922
rect -784 4888 -748 4922
rect -714 4888 -678 4922
rect -644 4888 -608 4922
rect -574 4888 -538 4922
rect -504 4888 -468 4922
rect -434 4888 -398 4922
rect -364 4888 -328 4922
rect -294 4888 -258 4922
rect -224 4888 -188 4922
rect -154 4888 -118 4922
rect -84 4888 -48 4922
rect -14 4918 102 4922
rect -14 4888 68 4918
rect -852 4884 68 4888
rect -852 4854 102 4884
rect -852 4820 -818 4854
rect -784 4820 -748 4854
rect -714 4820 -678 4854
rect -644 4820 -608 4854
rect -574 4820 -538 4854
rect -504 4820 -468 4854
rect -434 4820 -398 4854
rect -364 4820 -328 4854
rect -294 4820 -258 4854
rect -224 4820 -188 4854
rect -154 4820 -118 4854
rect -84 4820 -48 4854
rect -14 4850 102 4854
rect -14 4820 68 4850
rect -852 4816 68 4820
rect -852 4786 102 4816
rect -852 4752 -818 4786
rect -784 4752 -748 4786
rect -714 4752 -678 4786
rect -644 4752 -608 4786
rect -574 4752 -538 4786
rect -504 4752 -468 4786
rect -434 4752 -398 4786
rect -364 4752 -328 4786
rect -294 4752 -258 4786
rect -224 4752 -188 4786
rect -154 4752 -118 4786
rect -84 4752 -48 4786
rect -14 4782 102 4786
rect -14 4752 68 4782
rect -852 4748 68 4752
rect -852 4718 102 4748
rect -852 4684 -818 4718
rect -784 4684 -748 4718
rect -714 4684 -678 4718
rect -644 4684 -608 4718
rect -574 4684 -538 4718
rect -504 4684 -468 4718
rect -434 4684 -398 4718
rect -364 4684 -328 4718
rect -294 4684 -258 4718
rect -224 4684 -188 4718
rect -154 4684 -118 4718
rect -84 4684 -48 4718
rect -14 4714 102 4718
rect -14 4684 68 4714
rect -852 4680 68 4684
rect -852 4650 102 4680
rect -852 4616 -818 4650
rect -784 4616 -748 4650
rect -714 4616 -678 4650
rect -644 4616 -608 4650
rect -574 4616 -538 4650
rect -504 4616 -468 4650
rect -434 4616 -398 4650
rect -364 4616 -328 4650
rect -294 4616 -258 4650
rect -224 4616 -188 4650
rect -154 4616 -118 4650
rect -84 4616 -48 4650
rect -14 4646 102 4650
rect -14 4616 68 4646
rect -852 4612 68 4616
rect -852 4582 102 4612
rect -852 4548 -818 4582
rect -784 4548 -748 4582
rect -714 4548 -678 4582
rect -644 4548 -608 4582
rect -574 4548 -538 4582
rect -504 4548 -468 4582
rect -434 4548 -398 4582
rect -364 4548 -328 4582
rect -294 4548 -258 4582
rect -224 4548 -188 4582
rect -154 4548 -118 4582
rect -84 4548 -48 4582
rect -14 4578 102 4582
rect -14 4548 68 4578
rect -852 4544 68 4548
rect -852 4514 102 4544
rect -852 4480 -818 4514
rect -784 4480 -748 4514
rect -714 4480 -678 4514
rect -644 4480 -608 4514
rect -574 4480 -538 4514
rect -504 4480 -468 4514
rect -434 4480 -398 4514
rect -364 4480 -328 4514
rect -294 4480 -258 4514
rect -224 4480 -188 4514
rect -154 4480 -118 4514
rect -84 4480 -48 4514
rect -14 4510 102 4514
rect -14 4480 68 4510
rect -852 4476 68 4480
rect -852 4446 102 4476
rect -852 4412 -818 4446
rect -784 4412 -748 4446
rect -714 4412 -678 4446
rect -644 4412 -608 4446
rect -574 4412 -538 4446
rect -504 4412 -468 4446
rect -434 4412 -398 4446
rect -364 4412 -328 4446
rect -294 4412 -258 4446
rect -224 4412 -188 4446
rect -154 4412 -118 4446
rect -84 4412 -48 4446
rect -14 4442 102 4446
rect -14 4412 68 4442
rect -852 4408 68 4412
rect -852 4378 102 4408
rect -852 4344 -818 4378
rect -784 4344 -748 4378
rect -714 4344 -678 4378
rect -644 4344 -608 4378
rect -574 4344 -538 4378
rect -504 4344 -468 4378
rect -434 4344 -398 4378
rect -364 4344 -328 4378
rect -294 4344 -258 4378
rect -224 4344 -188 4378
rect -154 4344 -118 4378
rect -84 4344 -48 4378
rect -14 4374 102 4378
rect -14 4344 68 4374
rect -852 4340 68 4344
rect -852 4310 102 4340
rect -852 4276 -818 4310
rect -784 4276 -748 4310
rect -714 4276 -678 4310
rect -644 4276 -608 4310
rect -574 4276 -538 4310
rect -504 4276 -468 4310
rect -434 4276 -398 4310
rect -364 4276 -328 4310
rect -294 4276 -258 4310
rect -224 4276 -188 4310
rect -154 4276 -118 4310
rect -84 4276 -48 4310
rect -14 4306 102 4310
rect -14 4276 68 4306
rect -852 4272 68 4276
rect -852 4242 102 4272
rect -852 4208 -818 4242
rect -784 4208 -748 4242
rect -714 4208 -678 4242
rect -644 4208 -608 4242
rect -574 4208 -538 4242
rect -504 4208 -468 4242
rect -434 4208 -398 4242
rect -364 4208 -328 4242
rect -294 4208 -258 4242
rect -224 4208 -188 4242
rect -154 4208 -118 4242
rect -84 4208 -48 4242
rect -14 4238 102 4242
rect -14 4208 68 4238
rect -852 4204 68 4208
rect -852 4174 102 4204
rect -852 4140 -818 4174
rect -784 4140 -748 4174
rect -714 4140 -678 4174
rect -644 4140 -608 4174
rect -574 4140 -538 4174
rect -504 4140 -468 4174
rect -434 4140 -398 4174
rect -364 4140 -328 4174
rect -294 4140 -258 4174
rect -224 4140 -188 4174
rect -154 4140 -118 4174
rect -84 4140 -48 4174
rect -14 4170 102 4174
rect -14 4140 68 4170
rect -852 4136 68 4140
rect -852 4106 102 4136
rect -852 4072 -818 4106
rect -784 4072 -748 4106
rect -714 4072 -678 4106
rect -644 4072 -608 4106
rect -574 4072 -538 4106
rect -504 4072 -468 4106
rect -434 4072 -398 4106
rect -364 4072 -328 4106
rect -294 4072 -258 4106
rect -224 4072 -188 4106
rect -154 4072 -118 4106
rect -84 4072 -48 4106
rect -14 4102 102 4106
rect -14 4072 68 4102
rect -852 4068 68 4072
rect -852 4038 102 4068
rect -852 4004 -818 4038
rect -784 4004 -748 4038
rect -714 4004 -678 4038
rect -644 4004 -608 4038
rect -574 4004 -538 4038
rect -504 4004 -468 4038
rect -434 4004 -398 4038
rect -364 4004 -328 4038
rect -294 4004 -258 4038
rect -224 4004 -188 4038
rect -154 4004 -118 4038
rect -84 4004 -48 4038
rect -14 4034 102 4038
rect -14 4004 68 4034
rect -852 4000 68 4004
rect -852 3970 102 4000
rect -852 3936 -818 3970
rect -784 3936 -748 3970
rect -714 3936 -678 3970
rect -644 3936 -608 3970
rect -574 3936 -538 3970
rect -504 3936 -468 3970
rect -434 3936 -398 3970
rect -364 3936 -328 3970
rect -294 3936 -258 3970
rect -224 3936 -188 3970
rect -154 3936 -118 3970
rect -84 3936 -48 3970
rect -14 3966 102 3970
rect -14 3936 68 3966
rect -852 3932 68 3936
rect -852 3902 102 3932
rect -852 3868 -818 3902
rect -784 3868 -748 3902
rect -714 3868 -678 3902
rect -644 3868 -608 3902
rect -574 3868 -538 3902
rect -504 3868 -468 3902
rect -434 3868 -398 3902
rect -364 3868 -328 3902
rect -294 3868 -258 3902
rect -224 3868 -188 3902
rect -154 3868 -118 3902
rect -84 3868 -48 3902
rect -14 3898 102 3902
rect -14 3868 68 3898
rect -852 3864 68 3868
rect -852 3834 102 3864
rect -852 3800 -818 3834
rect -784 3800 -748 3834
rect -714 3800 -678 3834
rect -644 3800 -608 3834
rect -574 3800 -538 3834
rect -504 3800 -468 3834
rect -434 3800 -398 3834
rect -364 3800 -328 3834
rect -294 3800 -258 3834
rect -224 3800 -188 3834
rect -154 3800 -118 3834
rect -84 3800 -48 3834
rect -14 3830 102 3834
rect -14 3800 68 3830
rect -852 3796 68 3800
rect -852 3766 102 3796
rect -852 3732 -818 3766
rect -784 3732 -748 3766
rect -714 3732 -678 3766
rect -644 3732 -608 3766
rect -574 3732 -538 3766
rect -504 3732 -468 3766
rect -434 3732 -398 3766
rect -364 3732 -328 3766
rect -294 3732 -258 3766
rect -224 3732 -188 3766
rect -154 3732 -118 3766
rect -84 3732 -48 3766
rect -14 3762 102 3766
rect -14 3732 68 3762
rect -852 3728 68 3732
rect -852 3698 102 3728
rect -852 3664 -818 3698
rect -784 3664 -748 3698
rect -714 3664 -678 3698
rect -644 3664 -608 3698
rect -574 3664 -538 3698
rect -504 3664 -468 3698
rect -434 3664 -398 3698
rect -364 3664 -328 3698
rect -294 3664 -258 3698
rect -224 3664 -188 3698
rect -154 3664 -118 3698
rect -84 3664 -48 3698
rect -14 3694 102 3698
rect -14 3664 68 3694
rect -852 3660 68 3664
rect -852 3630 102 3660
rect -852 3596 -818 3630
rect -784 3596 -748 3630
rect -714 3596 -678 3630
rect -644 3596 -608 3630
rect -574 3596 -538 3630
rect -504 3596 -468 3630
rect -434 3596 -398 3630
rect -364 3596 -328 3630
rect -294 3596 -258 3630
rect -224 3596 -188 3630
rect -154 3596 -118 3630
rect -84 3596 -48 3630
rect -14 3626 102 3630
rect -14 3596 68 3626
rect -852 3592 68 3596
rect -852 3562 102 3592
rect -852 3528 -818 3562
rect -784 3528 -748 3562
rect -714 3528 -678 3562
rect -644 3528 -608 3562
rect -574 3528 -538 3562
rect -504 3528 -468 3562
rect -434 3528 -398 3562
rect -364 3528 -328 3562
rect -294 3528 -258 3562
rect -224 3528 -188 3562
rect -154 3528 -118 3562
rect -84 3528 -48 3562
rect -14 3558 102 3562
rect -14 3528 68 3558
rect -852 3524 68 3528
rect -852 3494 102 3524
rect -852 3460 -818 3494
rect -784 3460 -748 3494
rect -714 3460 -678 3494
rect -644 3460 -608 3494
rect -574 3460 -538 3494
rect -504 3460 -468 3494
rect -434 3460 -398 3494
rect -364 3460 -328 3494
rect -294 3460 -258 3494
rect -224 3460 -188 3494
rect -154 3460 -118 3494
rect -84 3460 -48 3494
rect -14 3490 102 3494
rect -14 3460 68 3490
rect -852 3456 68 3460
rect -852 3426 102 3456
rect -852 3392 -818 3426
rect -784 3392 -748 3426
rect -714 3392 -678 3426
rect -644 3392 -608 3426
rect -574 3392 -538 3426
rect -504 3392 -468 3426
rect -434 3392 -398 3426
rect -364 3392 -328 3426
rect -294 3392 -258 3426
rect -224 3392 -188 3426
rect -154 3392 -118 3426
rect -84 3392 -48 3426
rect -14 3422 102 3426
rect -14 3392 68 3422
rect -852 3388 68 3392
rect -852 3358 102 3388
rect -852 3324 -818 3358
rect -784 3324 -748 3358
rect -714 3324 -678 3358
rect -644 3324 -608 3358
rect -574 3324 -538 3358
rect -504 3324 -468 3358
rect -434 3324 -398 3358
rect -364 3324 -328 3358
rect -294 3324 -258 3358
rect -224 3324 -188 3358
rect -154 3324 -118 3358
rect -84 3324 -48 3358
rect -14 3354 102 3358
rect -14 3324 68 3354
rect -852 3320 68 3324
rect -852 3290 102 3320
rect -852 3256 -818 3290
rect -784 3256 -748 3290
rect -714 3256 -678 3290
rect -644 3256 -608 3290
rect -574 3256 -538 3290
rect -504 3256 -468 3290
rect -434 3256 -398 3290
rect -364 3256 -328 3290
rect -294 3256 -258 3290
rect -224 3256 -188 3290
rect -154 3256 -118 3290
rect -84 3256 -48 3290
rect -14 3286 102 3290
rect -14 3256 68 3286
rect -852 3252 68 3256
rect -852 3222 102 3252
rect -852 3188 -818 3222
rect -784 3188 -748 3222
rect -714 3188 -678 3222
rect -644 3188 -608 3222
rect -574 3188 -538 3222
rect -504 3188 -468 3222
rect -434 3188 -398 3222
rect -364 3188 -328 3222
rect -294 3188 -258 3222
rect -224 3188 -188 3222
rect -154 3188 -118 3222
rect -84 3188 -48 3222
rect -14 3218 102 3222
rect -14 3188 68 3218
rect -852 3184 68 3188
rect -852 3154 102 3184
rect -852 3120 -818 3154
rect -784 3120 -748 3154
rect -714 3120 -678 3154
rect -644 3120 -608 3154
rect -574 3120 -538 3154
rect -504 3120 -468 3154
rect -434 3120 -398 3154
rect -364 3120 -328 3154
rect -294 3120 -258 3154
rect -224 3120 -188 3154
rect -154 3120 -118 3154
rect -84 3120 -48 3154
rect -14 3150 102 3154
rect -14 3120 68 3150
rect -852 3116 68 3120
rect -852 3086 102 3116
rect -852 3052 -818 3086
rect -784 3052 -748 3086
rect -714 3052 -678 3086
rect -644 3052 -608 3086
rect -574 3052 -538 3086
rect -504 3052 -468 3086
rect -434 3052 -398 3086
rect -364 3052 -328 3086
rect -294 3052 -258 3086
rect -224 3052 -188 3086
rect -154 3052 -118 3086
rect -84 3052 -48 3086
rect -14 3082 102 3086
rect -14 3052 68 3082
rect -852 3048 68 3052
rect -852 3018 102 3048
rect -852 2984 -818 3018
rect -784 2984 -748 3018
rect -714 2984 -678 3018
rect -644 2984 -608 3018
rect -574 2984 -538 3018
rect -504 2984 -468 3018
rect -434 2984 -398 3018
rect -364 2984 -328 3018
rect -294 2984 -258 3018
rect -224 2984 -188 3018
rect -154 2984 -118 3018
rect -84 2984 -48 3018
rect -14 3014 102 3018
rect -14 2984 68 3014
rect -852 2980 68 2984
rect -852 2950 102 2980
rect -852 2916 -818 2950
rect -784 2916 -748 2950
rect -714 2916 -678 2950
rect -644 2916 -608 2950
rect -574 2916 -538 2950
rect -504 2916 -468 2950
rect -434 2916 -398 2950
rect -364 2916 -328 2950
rect -294 2916 -258 2950
rect -224 2916 -188 2950
rect -154 2916 -118 2950
rect -84 2916 -48 2950
rect -14 2946 102 2950
rect -14 2916 68 2946
rect -852 2912 68 2916
rect -852 2882 102 2912
rect -852 2848 -818 2882
rect -784 2848 -748 2882
rect -714 2848 -678 2882
rect -644 2848 -608 2882
rect -574 2848 -538 2882
rect -504 2848 -468 2882
rect -434 2848 -398 2882
rect -364 2848 -328 2882
rect -294 2848 -258 2882
rect -224 2848 -188 2882
rect -154 2848 -118 2882
rect -84 2848 -48 2882
rect -14 2878 102 2882
rect -14 2848 68 2878
rect -852 2844 68 2848
rect -852 2814 102 2844
rect -852 2780 -818 2814
rect -784 2780 -748 2814
rect -714 2780 -678 2814
rect -644 2780 -608 2814
rect -574 2780 -538 2814
rect -504 2780 -468 2814
rect -434 2780 -398 2814
rect -364 2780 -328 2814
rect -294 2780 -258 2814
rect -224 2780 -188 2814
rect -154 2780 -118 2814
rect -84 2780 -48 2814
rect -14 2810 102 2814
rect -14 2780 68 2810
rect -852 2776 68 2780
rect -852 2746 102 2776
rect -852 2712 -818 2746
rect -784 2712 -748 2746
rect -714 2712 -678 2746
rect -644 2712 -608 2746
rect -574 2712 -538 2746
rect -504 2712 -468 2746
rect -434 2712 -398 2746
rect -364 2712 -328 2746
rect -294 2712 -258 2746
rect -224 2712 -188 2746
rect -154 2712 -118 2746
rect -84 2712 -48 2746
rect -14 2742 102 2746
rect -14 2712 68 2742
rect -852 2708 68 2712
rect -852 2678 102 2708
rect -852 2644 -818 2678
rect -784 2644 -748 2678
rect -714 2644 -678 2678
rect -644 2644 -608 2678
rect -574 2644 -538 2678
rect -504 2644 -468 2678
rect -434 2644 -398 2678
rect -364 2644 -328 2678
rect -294 2644 -258 2678
rect -224 2644 -188 2678
rect -154 2644 -118 2678
rect -84 2644 -48 2678
rect -14 2674 102 2678
rect -14 2644 68 2674
rect -852 2640 68 2644
rect -852 2610 102 2640
rect -852 2576 -818 2610
rect -784 2576 -748 2610
rect -714 2576 -678 2610
rect -644 2576 -608 2610
rect -574 2576 -538 2610
rect -504 2576 -468 2610
rect -434 2576 -398 2610
rect -364 2576 -328 2610
rect -294 2576 -258 2610
rect -224 2576 -188 2610
rect -154 2576 -118 2610
rect -84 2576 -48 2610
rect -14 2606 102 2610
rect -14 2576 68 2606
rect -852 2572 68 2576
rect -852 2542 102 2572
rect -852 2508 -818 2542
rect -784 2508 -748 2542
rect -714 2508 -678 2542
rect -644 2508 -608 2542
rect -574 2508 -538 2542
rect -504 2508 -468 2542
rect -434 2508 -398 2542
rect -364 2508 -328 2542
rect -294 2508 -258 2542
rect -224 2508 -188 2542
rect -154 2508 -118 2542
rect -84 2508 -48 2542
rect -14 2538 102 2542
rect -14 2508 68 2538
rect -852 2504 68 2508
rect -852 2473 102 2504
rect -852 2439 -818 2473
rect -784 2439 -748 2473
rect -714 2439 -678 2473
rect -644 2439 -608 2473
rect -574 2439 -538 2473
rect -504 2439 -468 2473
rect -434 2439 -398 2473
rect -364 2439 -328 2473
rect -294 2439 -258 2473
rect -224 2439 -188 2473
rect -154 2439 -118 2473
rect -84 2439 -48 2473
rect -14 2470 102 2473
rect -14 2439 68 2470
rect -852 2436 68 2439
rect -852 2404 102 2436
rect -852 2370 -818 2404
rect -784 2370 -748 2404
rect -714 2370 -678 2404
rect -644 2370 -608 2404
rect -574 2370 -538 2404
rect -504 2370 -468 2404
rect -434 2370 -398 2404
rect -364 2370 -328 2404
rect -294 2370 -258 2404
rect -224 2370 -188 2404
rect -154 2370 -118 2404
rect -84 2370 -48 2404
rect -14 2402 102 2404
rect -14 2370 68 2402
rect -852 2368 68 2370
rect -852 2335 102 2368
rect -852 2301 -818 2335
rect -784 2301 -748 2335
rect -714 2301 -678 2335
rect -644 2301 -608 2335
rect -574 2301 -538 2335
rect -504 2301 -468 2335
rect -434 2301 -398 2335
rect -364 2301 -328 2335
rect -294 2301 -258 2335
rect -224 2301 -188 2335
rect -154 2301 -118 2335
rect -84 2301 -48 2335
rect -14 2334 102 2335
rect -14 2301 68 2334
rect -852 2300 68 2301
rect -852 2266 102 2300
rect -852 2232 -818 2266
rect -784 2232 -748 2266
rect -714 2232 -678 2266
rect -644 2232 -608 2266
rect -574 2232 -538 2266
rect -504 2232 -468 2266
rect -434 2232 -398 2266
rect -364 2232 -328 2266
rect -294 2232 -258 2266
rect -224 2232 -188 2266
rect -154 2232 -118 2266
rect -84 2232 -48 2266
rect -14 2232 68 2266
rect -852 2198 102 2232
rect -852 2197 68 2198
rect -852 2163 -818 2197
rect -784 2163 -748 2197
rect -714 2163 -678 2197
rect -644 2163 -608 2197
rect -574 2163 -538 2197
rect -504 2163 -468 2197
rect -434 2163 -398 2197
rect -364 2163 -328 2197
rect -294 2163 -258 2197
rect -224 2163 -188 2197
rect -154 2163 -118 2197
rect -84 2163 -48 2197
rect -14 2164 68 2197
rect -14 2163 102 2164
rect -852 2130 102 2163
rect -852 2128 68 2130
rect -852 2094 -818 2128
rect -784 2094 -748 2128
rect -714 2094 -678 2128
rect -644 2094 -608 2128
rect -574 2094 -538 2128
rect -504 2094 -468 2128
rect -434 2094 -398 2128
rect -364 2094 -328 2128
rect -294 2094 -258 2128
rect -224 2094 -188 2128
rect -154 2094 -118 2128
rect -84 2094 -48 2128
rect -14 2096 68 2128
rect -14 2094 102 2096
rect -852 2062 102 2094
rect -852 2059 68 2062
rect -852 2025 -818 2059
rect -784 2025 -748 2059
rect -714 2025 -678 2059
rect -644 2025 -608 2059
rect -574 2025 -538 2059
rect -504 2025 -468 2059
rect -434 2025 -398 2059
rect -364 2025 -328 2059
rect -294 2025 -258 2059
rect -224 2025 -188 2059
rect -154 2025 -118 2059
rect -84 2025 -48 2059
rect -14 2028 68 2059
rect -14 2025 102 2028
rect -852 1994 102 2025
rect -852 1990 68 1994
rect -852 1956 -818 1990
rect -784 1956 -748 1990
rect -714 1956 -678 1990
rect -644 1956 -608 1990
rect -574 1956 -538 1990
rect -504 1956 -468 1990
rect -434 1956 -398 1990
rect -364 1956 -328 1990
rect -294 1956 -258 1990
rect -224 1956 -188 1990
rect -154 1956 -118 1990
rect -84 1956 -48 1990
rect -14 1960 68 1990
rect -14 1956 102 1960
rect -852 1926 102 1956
rect -852 1921 68 1926
rect -852 1887 -818 1921
rect -784 1887 -748 1921
rect -714 1887 -678 1921
rect -644 1887 -608 1921
rect -574 1887 -538 1921
rect -504 1887 -468 1921
rect -434 1887 -398 1921
rect -364 1887 -328 1921
rect -294 1887 -258 1921
rect -224 1887 -188 1921
rect -154 1887 -118 1921
rect -84 1887 -48 1921
rect -14 1892 68 1921
rect -14 1887 102 1892
rect -852 1858 102 1887
rect -852 1852 68 1858
rect -852 1818 -818 1852
rect -784 1818 -748 1852
rect -714 1818 -678 1852
rect -644 1818 -608 1852
rect -574 1818 -538 1852
rect -504 1818 -468 1852
rect -434 1818 -398 1852
rect -364 1818 -328 1852
rect -294 1818 -258 1852
rect -224 1818 -188 1852
rect -154 1818 -118 1852
rect -84 1818 -48 1852
rect -14 1824 68 1852
rect -14 1818 102 1824
rect -852 1790 102 1818
rect -852 1783 68 1790
rect -852 1749 -818 1783
rect -784 1749 -748 1783
rect -714 1749 -678 1783
rect -644 1749 -608 1783
rect -574 1749 -538 1783
rect -504 1749 -468 1783
rect -434 1749 -398 1783
rect -364 1749 -328 1783
rect -294 1749 -258 1783
rect -224 1749 -188 1783
rect -154 1749 -118 1783
rect -84 1749 -48 1783
rect -14 1756 68 1783
rect -14 1749 102 1756
rect -852 1722 102 1749
rect -852 1714 68 1722
rect -852 1680 -818 1714
rect -784 1680 -748 1714
rect -714 1680 -678 1714
rect -644 1680 -608 1714
rect -574 1680 -538 1714
rect -504 1680 -468 1714
rect -434 1680 -398 1714
rect -364 1680 -328 1714
rect -294 1680 -258 1714
rect -224 1680 -188 1714
rect -154 1680 -118 1714
rect -84 1680 -48 1714
rect -14 1688 68 1714
rect -14 1680 102 1688
rect -852 1654 102 1680
rect -852 1645 68 1654
rect -852 1611 -818 1645
rect -784 1611 -748 1645
rect -714 1611 -678 1645
rect -644 1611 -608 1645
rect -574 1611 -538 1645
rect -504 1611 -468 1645
rect -434 1611 -398 1645
rect -364 1611 -328 1645
rect -294 1611 -258 1645
rect -224 1611 -188 1645
rect -154 1611 -118 1645
rect -84 1611 -48 1645
rect -14 1620 68 1645
rect -14 1611 102 1620
rect -852 1586 102 1611
rect -852 1576 68 1586
rect -852 1542 -818 1576
rect -784 1542 -748 1576
rect -714 1542 -678 1576
rect -644 1542 -608 1576
rect -574 1542 -538 1576
rect -504 1542 -468 1576
rect -434 1542 -398 1576
rect -364 1542 -328 1576
rect -294 1542 -258 1576
rect -224 1542 -188 1576
rect -154 1542 -118 1576
rect -84 1542 -48 1576
rect -14 1552 68 1576
rect -14 1542 102 1552
rect -852 1518 102 1542
rect -852 1507 68 1518
rect -852 1473 -818 1507
rect -784 1473 -748 1507
rect -714 1473 -678 1507
rect -644 1473 -608 1507
rect -574 1473 -538 1507
rect -504 1473 -468 1507
rect -434 1473 -398 1507
rect -364 1473 -328 1507
rect -294 1473 -258 1507
rect -224 1473 -188 1507
rect -154 1473 -118 1507
rect -84 1473 -48 1507
rect -14 1484 68 1507
rect -14 1473 102 1484
rect -852 1450 102 1473
rect -852 1438 68 1450
rect -852 1404 -818 1438
rect -784 1404 -748 1438
rect -714 1404 -678 1438
rect -644 1404 -608 1438
rect -574 1404 -538 1438
rect -504 1404 -468 1438
rect -434 1404 -398 1438
rect -364 1404 -328 1438
rect -294 1404 -258 1438
rect -224 1404 -188 1438
rect -154 1404 -118 1438
rect -84 1404 -48 1438
rect -14 1416 68 1438
rect -14 1404 102 1416
rect -852 1381 102 1404
rect -852 1369 68 1381
rect -852 1335 -818 1369
rect -784 1335 -748 1369
rect -714 1335 -678 1369
rect -644 1335 -608 1369
rect -574 1335 -538 1369
rect -504 1335 -468 1369
rect -434 1335 -398 1369
rect -364 1335 -328 1369
rect -294 1335 -258 1369
rect -224 1335 -188 1369
rect -154 1335 -118 1369
rect -84 1335 -48 1369
rect -14 1347 68 1369
rect -14 1335 102 1347
rect -852 1312 102 1335
rect -852 1300 68 1312
rect -852 1266 -818 1300
rect -784 1266 -748 1300
rect -714 1266 -678 1300
rect -644 1266 -608 1300
rect -574 1266 -538 1300
rect -504 1266 -468 1300
rect -434 1266 -398 1300
rect -364 1266 -328 1300
rect -294 1266 -258 1300
rect -224 1266 -188 1300
rect -154 1266 -118 1300
rect -84 1266 -48 1300
rect -14 1278 68 1300
rect -14 1266 102 1278
rect -852 1243 102 1266
rect -852 1231 68 1243
rect -852 1197 -818 1231
rect -784 1197 -748 1231
rect -714 1197 -678 1231
rect -644 1197 -608 1231
rect -574 1197 -538 1231
rect -504 1197 -468 1231
rect -434 1197 -398 1231
rect -364 1197 -328 1231
rect -294 1197 -258 1231
rect -224 1197 -188 1231
rect -154 1197 -118 1231
rect -84 1197 -48 1231
rect -14 1209 68 1231
rect -14 1197 102 1209
rect -852 1174 102 1197
rect -852 1162 68 1174
rect -852 1128 -818 1162
rect -784 1128 -748 1162
rect -714 1128 -678 1162
rect -644 1128 -608 1162
rect -574 1128 -538 1162
rect -504 1128 -468 1162
rect -434 1128 -398 1162
rect -364 1128 -328 1162
rect -294 1128 -258 1162
rect -224 1128 -188 1162
rect -154 1128 -118 1162
rect -84 1128 -48 1162
rect -14 1140 68 1162
rect -14 1128 102 1140
rect -852 1105 102 1128
rect -852 1093 68 1105
rect -852 1059 -818 1093
rect -784 1059 -748 1093
rect -714 1059 -678 1093
rect -644 1059 -608 1093
rect -574 1059 -538 1093
rect -504 1059 -468 1093
rect -434 1059 -398 1093
rect -364 1059 -328 1093
rect -294 1059 -258 1093
rect -224 1059 -188 1093
rect -154 1059 -118 1093
rect -84 1059 -48 1093
rect -14 1071 68 1093
rect -14 1059 102 1071
rect -852 1036 102 1059
rect -852 1024 68 1036
rect -852 990 -818 1024
rect -784 990 -748 1024
rect -714 990 -678 1024
rect -644 990 -608 1024
rect -574 990 -538 1024
rect -504 990 -468 1024
rect -434 990 -398 1024
rect -364 990 -328 1024
rect -294 990 -258 1024
rect -224 990 -188 1024
rect -154 990 -118 1024
rect -84 990 -48 1024
rect -14 1002 68 1024
rect -14 990 102 1002
rect -852 967 102 990
rect -852 955 68 967
rect -852 921 -818 955
rect -784 921 -748 955
rect -714 921 -678 955
rect -644 921 -608 955
rect -574 921 -538 955
rect -504 921 -468 955
rect -434 921 -398 955
rect -364 921 -328 955
rect -294 921 -258 955
rect -224 921 -188 955
rect -154 921 -118 955
rect -84 921 -48 955
rect -14 933 68 955
rect -14 921 102 933
rect -852 898 102 921
rect -852 886 68 898
rect -852 852 -818 886
rect -784 852 -748 886
rect -714 852 -678 886
rect -644 852 -608 886
rect -574 852 -538 886
rect -504 852 -468 886
rect -434 852 -398 886
rect -364 852 -328 886
rect -294 852 -258 886
rect -224 852 -188 886
rect -154 852 -118 886
rect -84 852 -48 886
rect -14 864 68 886
rect -14 852 102 864
rect -852 829 102 852
rect -852 817 68 829
rect -852 783 -818 817
rect -784 783 -748 817
rect -714 783 -678 817
rect -644 783 -608 817
rect -574 783 -538 817
rect -504 783 -468 817
rect -434 783 -398 817
rect -364 783 -328 817
rect -294 783 -258 817
rect -224 783 -188 817
rect -154 783 -118 817
rect -84 783 -48 817
rect -14 795 68 817
rect -14 783 102 795
rect -852 760 102 783
rect -852 748 68 760
rect -852 714 -818 748
rect -784 714 -748 748
rect -714 714 -678 748
rect -644 714 -608 748
rect -574 714 -538 748
rect -504 714 -468 748
rect -434 714 -398 748
rect -364 714 -328 748
rect -294 714 -258 748
rect -224 714 -188 748
rect -154 714 -118 748
rect -84 714 -48 748
rect -14 726 68 748
rect -14 714 102 726
rect -852 691 102 714
rect -852 679 68 691
rect -852 645 -818 679
rect -784 645 -748 679
rect -714 645 -678 679
rect -644 645 -608 679
rect -574 645 -538 679
rect -504 645 -468 679
rect -434 645 -398 679
rect -364 645 -328 679
rect -294 645 -258 679
rect -224 645 -188 679
rect -154 645 -118 679
rect -84 645 -48 679
rect -14 657 68 679
rect -14 645 102 657
rect -852 622 102 645
rect -852 610 68 622
rect -852 576 -818 610
rect -784 576 -748 610
rect -714 576 -678 610
rect -644 576 -608 610
rect -574 576 -538 610
rect -504 576 -468 610
rect -434 576 -398 610
rect -364 576 -328 610
rect -294 576 -258 610
rect -224 576 -188 610
rect -154 576 -118 610
rect -84 576 -48 610
rect -14 588 68 610
rect -14 576 102 588
rect -852 553 102 576
rect -852 541 68 553
rect -852 507 -818 541
rect -784 507 -748 541
rect -714 507 -678 541
rect -644 507 -608 541
rect -574 507 -538 541
rect -504 507 -468 541
rect -434 507 -398 541
rect -364 507 -328 541
rect -294 507 -258 541
rect -224 507 -188 541
rect -154 507 -118 541
rect -84 507 -48 541
rect -14 519 68 541
rect -14 507 102 519
rect -852 484 102 507
rect -852 472 68 484
rect -852 438 -818 472
rect -784 438 -748 472
rect -714 438 -678 472
rect -644 438 -608 472
rect -574 438 -538 472
rect -504 438 -468 472
rect -434 438 -398 472
rect -364 438 -328 472
rect -294 438 -258 472
rect -224 438 -188 472
rect -154 438 -118 472
rect -84 438 -48 472
rect -14 450 68 472
rect -14 438 102 450
rect -852 415 102 438
rect -852 403 68 415
rect -852 369 -818 403
rect -784 369 -748 403
rect -714 369 -678 403
rect -644 369 -608 403
rect -574 369 -538 403
rect -504 369 -468 403
rect -434 369 -398 403
rect -364 369 -328 403
rect -294 369 -258 403
rect -224 369 -188 403
rect -154 369 -118 403
rect -84 369 -48 403
rect -14 381 68 403
rect -14 369 102 381
rect -852 346 102 369
rect -852 334 68 346
rect -852 300 -818 334
rect -784 300 -748 334
rect -714 300 -678 334
rect -644 300 -608 334
rect -574 300 -538 334
rect -504 300 -468 334
rect -434 300 -398 334
rect -364 300 -328 334
rect -294 300 -258 334
rect -224 300 -188 334
rect -154 300 -118 334
rect -84 300 -48 334
rect -14 312 68 334
rect -14 300 102 312
rect -852 277 102 300
rect -852 265 68 277
rect -852 231 -818 265
rect -784 231 -748 265
rect -714 231 -678 265
rect -644 231 -608 265
rect -574 231 -538 265
rect -504 231 -468 265
rect -434 231 -398 265
rect -364 231 -328 265
rect -294 231 -258 265
rect -224 231 -188 265
rect -154 231 -118 265
rect -84 231 -48 265
rect -14 243 68 265
rect -14 231 102 243
rect -852 208 102 231
rect -852 196 68 208
rect -852 162 -818 196
rect -784 162 -748 196
rect -714 162 -678 196
rect -644 162 -608 196
rect -574 162 -538 196
rect -504 162 -468 196
rect -434 162 -398 196
rect -364 162 -328 196
rect -294 162 -258 196
rect -224 162 -188 196
rect -154 162 -118 196
rect -84 162 -48 196
rect -14 174 68 196
rect -14 162 102 174
rect -852 127 102 162
rect -852 93 -818 127
rect -784 93 -748 127
rect -714 93 -678 127
rect -644 93 -608 127
rect -574 93 -538 127
rect -504 93 -468 127
rect -434 93 -398 127
rect -364 93 -328 127
rect -294 93 -258 127
rect -224 93 -188 127
rect -154 93 -118 127
rect -84 93 -48 127
rect -14 102 102 127
rect 848 102 882 4976
rect -14 93 92 102
rect -852 68 92 93
rect 126 68 161 102
rect 195 68 230 102
rect 264 68 300 102
rect 334 68 370 102
rect 404 68 440 102
rect 474 68 510 102
rect 544 68 580 102
rect 614 68 650 102
rect 684 68 720 102
rect 754 68 790 102
rect 824 68 882 102
rect -852 58 882 68
rect -852 24 -818 58
rect -784 24 -748 58
rect -714 24 -678 58
rect -644 24 -608 58
rect -574 24 -538 58
rect -504 24 -468 58
rect -434 24 -398 58
rect -364 24 -328 58
rect -294 24 -258 58
rect -224 24 -188 58
rect -154 24 -118 58
rect -84 24 -48 58
rect -14 34 882 58
rect -14 24 92 34
rect -852 0 92 24
rect 126 0 161 34
rect 195 0 230 34
rect 264 0 300 34
rect 334 0 370 34
rect 404 0 440 34
rect 474 0 510 34
rect 544 0 580 34
rect 614 0 650 34
rect 684 0 720 34
rect 754 0 790 34
rect 824 0 882 34
rect -852 -33 882 0
rect -852 -34 898 -33
rect -852 -68 -818 -34
rect -784 -68 -750 -34
rect -716 -68 -682 -34
rect -648 -68 -614 -34
rect -580 -68 -546 -34
rect -512 -68 -478 -34
rect -444 -68 -410 -34
rect -376 -68 -342 -34
rect -308 -68 -274 -34
rect -240 -68 -205 -34
rect -171 -68 -136 -34
rect -102 -68 -67 -34
rect -33 -68 2 -34
rect 36 -68 71 -34
rect 105 -68 140 -34
rect 174 -68 209 -34
rect 243 -68 278 -34
rect 312 -68 347 -34
rect 381 -68 416 -34
rect 450 -68 485 -34
rect 519 -68 554 -34
rect 588 -68 623 -34
rect 657 -68 692 -34
rect 726 -68 761 -34
rect 795 -68 830 -34
rect 864 -68 898 -34
rect -852 -105 898 -68
rect -852 -139 -818 -105
rect -784 -139 -750 -105
rect -716 -139 -682 -105
rect -648 -139 -614 -105
rect -580 -139 -546 -105
rect -512 -139 -478 -105
rect -444 -139 -410 -105
rect -376 -139 -342 -105
rect -308 -139 -274 -105
rect -240 -139 -205 -105
rect -171 -139 -136 -105
rect -102 -139 -67 -105
rect -33 -139 2 -105
rect 36 -139 71 -105
rect 105 -139 140 -105
rect 174 -139 209 -105
rect 243 -139 278 -105
rect 312 -139 347 -105
rect 381 -139 416 -105
rect 450 -139 485 -105
rect 519 -139 554 -105
rect 588 -139 623 -105
rect 657 -139 692 -105
rect 726 -139 761 -105
rect 795 -139 830 -105
rect 864 -139 898 -105
rect -852 -176 898 -139
rect -852 -210 -818 -176
rect -784 -210 -750 -176
rect -716 -210 -682 -176
rect -648 -210 -614 -176
rect -580 -210 -546 -176
rect -512 -210 -478 -176
rect -444 -210 -410 -176
rect -376 -210 -342 -176
rect -308 -210 -274 -176
rect -240 -210 -205 -176
rect -171 -210 -136 -176
rect -102 -210 -67 -176
rect -33 -210 2 -176
rect 36 -210 71 -176
rect 105 -210 140 -176
rect 174 -210 209 -176
rect 243 -210 278 -176
rect 312 -210 347 -176
rect 381 -210 416 -176
rect 450 -210 485 -176
rect 519 -210 554 -176
rect 588 -210 623 -176
rect 657 -210 692 -176
rect 726 -210 761 -176
rect 795 -210 830 -176
rect 864 -210 898 -176
rect -852 -247 898 -210
rect -852 -281 -818 -247
rect -784 -281 -750 -247
rect -716 -281 -682 -247
rect -648 -281 -614 -247
rect -580 -281 -546 -247
rect -512 -281 -478 -247
rect -444 -281 -410 -247
rect -376 -281 -342 -247
rect -308 -281 -274 -247
rect -240 -281 -205 -247
rect -171 -281 -136 -247
rect -102 -281 -67 -247
rect -33 -281 2 -247
rect 36 -281 71 -247
rect 105 -281 140 -247
rect 174 -281 209 -247
rect 243 -281 278 -247
rect 312 -281 347 -247
rect 381 -281 416 -247
rect 450 -281 485 -247
rect 519 -281 554 -247
rect 588 -281 623 -247
rect 657 -281 692 -247
rect 726 -281 761 -247
rect 795 -281 830 -247
rect 864 -281 898 -247
rect -852 -318 898 -281
rect -852 -352 -818 -318
rect -784 -352 -750 -318
rect -716 -352 -682 -318
rect -648 -352 -614 -318
rect -580 -352 -546 -318
rect -512 -352 -478 -318
rect -444 -352 -410 -318
rect -376 -352 -342 -318
rect -308 -352 -274 -318
rect -240 -352 -205 -318
rect -171 -352 -136 -318
rect -102 -352 -67 -318
rect -33 -352 2 -318
rect 36 -352 71 -318
rect 105 -352 140 -318
rect 174 -352 209 -318
rect 243 -352 278 -318
rect 312 -352 347 -318
rect 381 -352 416 -318
rect 450 -352 485 -318
rect 519 -352 554 -318
rect 588 -352 623 -318
rect 657 -352 692 -318
rect 726 -352 761 -318
rect 795 -352 830 -318
rect 864 -352 898 -318
rect -852 -353 898 -352
<< mvpsubdiffcont >>
rect 278 4788 312 4822
rect 391 4788 425 4822
rect 525 4788 559 4822
rect 662 4764 696 4798
rect 254 4694 288 4728
rect 254 4625 288 4659
rect 254 4556 288 4590
rect 254 4487 288 4521
rect 254 4418 288 4452
rect 254 4349 288 4383
rect 254 4280 288 4314
rect 254 4211 288 4245
rect 254 4142 288 4176
rect 254 4073 288 4107
rect 254 4004 288 4038
rect 254 3935 288 3969
rect 254 3866 288 3900
rect 254 3797 288 3831
rect 254 3728 288 3762
rect 662 4695 696 4729
rect 662 4626 696 4660
rect 662 4557 696 4591
rect 662 4488 696 4522
rect 662 4419 696 4453
rect 662 4350 696 4384
rect 662 4281 696 4315
rect 662 4212 696 4246
rect 662 4143 696 4177
rect 662 4074 696 4108
rect 662 4005 696 4039
rect 662 3936 696 3970
rect 662 3867 696 3901
rect 662 3798 696 3832
rect 662 3729 696 3763
rect 254 3659 288 3693
rect 254 3590 288 3624
rect 662 3660 696 3694
rect 254 3521 288 3555
rect 254 3452 288 3486
rect 254 3383 288 3417
rect 254 3314 288 3348
rect 254 3245 288 3279
rect 254 3176 288 3210
rect 254 3107 288 3141
rect 254 3038 288 3072
rect 254 2969 288 3003
rect 254 2900 288 2934
rect 254 2831 288 2865
rect 254 2762 288 2796
rect 254 2693 288 2727
rect 254 2624 288 2658
rect 662 3591 696 3625
rect 662 3522 696 3556
rect 662 3453 696 3487
rect 662 3384 696 3418
rect 662 3315 696 3349
rect 662 3246 696 3280
rect 662 3177 696 3211
rect 662 3108 696 3142
rect 662 3039 696 3073
rect 662 2970 696 3004
rect 662 2901 696 2935
rect 662 2832 696 2866
rect 662 2763 696 2797
rect 662 2694 696 2728
rect 662 2625 696 2659
rect 254 2555 288 2589
rect 254 2486 288 2520
rect 662 2556 696 2590
rect 662 2487 696 2521
rect 254 2417 288 2451
rect 254 2348 288 2382
rect 254 2279 288 2313
rect 254 2210 288 2244
rect 254 2141 288 2175
rect 254 2072 288 2106
rect 254 2003 288 2037
rect 254 1934 288 1968
rect 254 1865 288 1899
rect 254 1796 288 1830
rect 254 1727 288 1761
rect 254 1658 288 1692
rect 254 1589 288 1623
rect 254 1520 288 1554
rect 254 1451 288 1485
rect 662 2418 696 2452
rect 662 2349 696 2383
rect 662 2280 696 2314
rect 662 2211 696 2245
rect 662 2142 696 2176
rect 662 2073 696 2107
rect 662 2004 696 2038
rect 662 1935 696 1969
rect 662 1866 696 1900
rect 662 1797 696 1831
rect 662 1728 696 1762
rect 662 1659 696 1693
rect 662 1590 696 1624
rect 662 1521 696 1555
rect 254 1382 288 1416
rect 662 1452 696 1486
rect 662 1383 696 1417
rect 254 1313 288 1347
rect 254 1244 288 1278
rect 254 1175 288 1209
rect 254 1106 288 1140
rect 254 1037 288 1071
rect 254 968 288 1002
rect 254 899 288 933
rect 254 830 288 864
rect 254 761 288 795
rect 254 692 288 726
rect 254 623 288 657
rect 254 554 288 588
rect 254 485 288 519
rect 254 416 288 450
rect 254 347 288 381
rect 662 1314 696 1348
rect 662 1245 696 1279
rect 662 1176 696 1210
rect 662 1107 696 1141
rect 662 1038 696 1072
rect 662 969 696 1003
rect 662 900 696 934
rect 662 831 696 865
rect 662 762 696 796
rect 662 693 696 727
rect 662 624 696 658
rect 662 555 696 589
rect 662 486 696 520
rect 662 417 696 451
rect 662 348 696 382
rect 254 278 288 312
rect 352 254 386 288
rect 423 254 457 288
rect 494 254 528 288
rect 566 254 600 288
rect 638 254 672 288
<< mvnsubdiffcont >>
rect -828 14648 -794 14682
rect -759 14648 -725 14682
rect -690 14648 -656 14682
rect -621 14648 -587 14682
rect -552 14648 -518 14682
rect -483 14648 -449 14682
rect -414 14648 -380 14682
rect -345 14648 -311 14682
rect -276 14648 -242 14682
rect -207 14648 -173 14682
rect -138 14648 -104 14682
rect -69 14648 -35 14682
rect 0 14648 34 14682
rect 69 14648 103 14682
rect 138 14648 172 14682
rect 207 14648 241 14682
rect 276 14648 310 14682
rect 345 14648 379 14682
rect 414 14648 448 14682
rect 483 14648 517 14682
rect 552 14648 586 14682
rect 621 14648 655 14682
rect 690 14648 724 14682
rect 759 14648 793 14682
rect 828 14648 862 14682
rect -828 14576 -794 14610
rect -759 14576 -725 14610
rect -690 14576 -656 14610
rect -621 14576 -587 14610
rect -552 14576 -518 14610
rect -483 14576 -449 14610
rect -414 14576 -380 14610
rect -345 14576 -311 14610
rect -276 14576 -242 14610
rect -207 14576 -173 14610
rect -138 14576 -104 14610
rect -69 14576 -35 14610
rect 0 14576 34 14610
rect 69 14576 103 14610
rect 138 14576 172 14610
rect 207 14576 241 14610
rect 276 14576 310 14610
rect 345 14576 379 14610
rect 414 14576 448 14610
rect 483 14576 517 14610
rect 552 14576 586 14610
rect 621 14576 655 14610
rect 690 14576 724 14610
rect 759 14576 793 14610
rect 828 14576 862 14610
rect -828 14504 -794 14538
rect -759 14504 -725 14538
rect -690 14504 -656 14538
rect -621 14504 -587 14538
rect -552 14504 -518 14538
rect -483 14504 -449 14538
rect -414 14504 -380 14538
rect -345 14504 -311 14538
rect -276 14504 -242 14538
rect -207 14504 -173 14538
rect -138 14504 -104 14538
rect -69 14504 -35 14538
rect 0 14504 34 14538
rect 69 14504 103 14538
rect 138 14504 172 14538
rect 207 14504 241 14538
rect 276 14504 310 14538
rect 345 14504 379 14538
rect 414 14504 448 14538
rect 483 14504 517 14538
rect 552 14504 586 14538
rect 621 14504 655 14538
rect 690 14504 724 14538
rect 759 14504 793 14538
rect 828 14504 862 14538
rect -828 14432 -794 14466
rect -759 14432 -725 14466
rect -690 14432 -656 14466
rect -621 14432 -587 14466
rect -552 14432 -518 14466
rect -483 14432 -449 14466
rect -414 14432 -380 14466
rect -345 14432 -311 14466
rect -276 14432 -242 14466
rect -207 14432 -173 14466
rect -138 14432 -104 14466
rect -69 14432 -35 14466
rect 0 14432 34 14466
rect 69 14432 103 14466
rect 138 14432 172 14466
rect 207 14432 241 14466
rect 276 14432 310 14466
rect 345 14432 379 14466
rect 414 14432 448 14466
rect 483 14432 517 14466
rect 552 14432 586 14466
rect 621 14432 655 14466
rect 690 14432 724 14466
rect 759 14432 793 14466
rect 828 14432 862 14466
rect -828 14360 -794 14394
rect -759 14360 -725 14394
rect -690 14360 -656 14394
rect -621 14360 -587 14394
rect -552 14360 -518 14394
rect -483 14360 -449 14394
rect -414 14360 -380 14394
rect -345 14360 -311 14394
rect -276 14360 -242 14394
rect -207 14360 -173 14394
rect -138 14360 -104 14394
rect -69 14360 -35 14394
rect 0 14360 34 14394
rect 69 14360 103 14394
rect 138 14360 172 14394
rect 207 14360 241 14394
rect 276 14360 310 14394
rect 345 14360 379 14394
rect 414 14360 448 14394
rect 483 14360 517 14394
rect 552 14360 586 14394
rect 621 14360 655 14394
rect 690 14360 724 14394
rect 759 14360 793 14394
rect 828 14360 862 14394
rect -828 14288 -794 14322
rect -759 14288 -725 14322
rect -690 14288 -656 14322
rect -621 14288 -587 14322
rect -552 14288 -518 14322
rect -483 14288 -449 14322
rect -414 14288 -380 14322
rect -345 14288 -311 14322
rect -276 14288 -242 14322
rect -207 14288 -173 14322
rect -138 14288 -104 14322
rect -69 14288 -35 14322
rect 0 14288 34 14322
rect 69 14288 103 14322
rect 138 14288 172 14322
rect 207 14288 241 14322
rect 276 14288 310 14322
rect 345 14288 379 14322
rect 414 14288 448 14322
rect 483 14288 517 14322
rect 552 14288 586 14322
rect 621 14288 655 14322
rect 690 14288 724 14322
rect 759 14288 793 14322
rect 828 14288 862 14322
rect -828 14216 -794 14250
rect -759 14216 -725 14250
rect -690 14216 -656 14250
rect -621 14216 -587 14250
rect -552 14216 -518 14250
rect -483 14216 -449 14250
rect -414 14216 -380 14250
rect -345 14216 -311 14250
rect -276 14216 -242 14250
rect -207 14216 -173 14250
rect -138 14216 -104 14250
rect -69 14216 -35 14250
rect 0 14216 34 14250
rect 69 14216 103 14250
rect 138 14216 172 14250
rect 207 14216 241 14250
rect 276 14216 310 14250
rect 345 14216 379 14250
rect 414 14216 448 14250
rect 483 14216 517 14250
rect 552 14216 586 14250
rect 621 14216 655 14250
rect 690 14216 724 14250
rect 759 14216 793 14250
rect 828 14216 862 14250
rect -828 14144 -794 14178
rect -759 14144 -725 14178
rect -690 14144 -656 14178
rect -621 14144 -587 14178
rect -552 14144 -518 14178
rect -483 14144 -449 14178
rect -414 14144 -380 14178
rect -345 14144 -311 14178
rect -276 14144 -242 14178
rect -207 14144 -173 14178
rect -138 14144 -104 14178
rect -69 14144 -35 14178
rect 0 14144 34 14178
rect 69 14144 103 14178
rect 138 14144 172 14178
rect 207 14144 241 14178
rect 276 14144 310 14178
rect 345 14144 379 14178
rect 414 14144 448 14178
rect 483 14144 517 14178
rect 552 14144 586 14178
rect 621 14144 655 14178
rect 690 14144 724 14178
rect 759 14144 793 14178
rect 828 14144 862 14178
rect -828 14072 -794 14106
rect -759 14072 -725 14106
rect -690 14072 -656 14106
rect -621 14072 -587 14106
rect -552 14072 -518 14106
rect -483 14072 -449 14106
rect -414 14072 -380 14106
rect -345 14072 -311 14106
rect -276 14072 -242 14106
rect -207 14072 -173 14106
rect -138 14072 -104 14106
rect -69 14072 -35 14106
rect 0 14072 34 14106
rect 69 14072 103 14106
rect 138 14072 172 14106
rect 207 14072 241 14106
rect 276 14072 310 14106
rect 345 14072 379 14106
rect 414 14072 448 14106
rect 483 14072 517 14106
rect 552 14072 586 14106
rect 621 14072 655 14106
rect 690 14072 724 14106
rect 759 14072 793 14106
rect 828 14072 862 14106
rect -828 14000 -794 14034
rect -759 14000 -725 14034
rect -690 14000 -656 14034
rect -621 14000 -587 14034
rect -552 14000 -518 14034
rect -483 14000 -449 14034
rect -414 14000 -380 14034
rect -345 14000 -311 14034
rect -276 14000 -242 14034
rect -207 14000 -173 14034
rect -138 14000 -104 14034
rect -69 14000 -35 14034
rect 0 14000 34 14034
rect 69 14000 103 14034
rect 138 14000 172 14034
rect 207 14000 241 14034
rect 276 14000 310 14034
rect 345 14000 379 14034
rect 414 14000 448 14034
rect 483 14000 517 14034
rect 552 14000 586 14034
rect 621 14000 655 14034
rect 690 14000 724 14034
rect 759 14000 793 14034
rect 828 14000 862 14034
rect -818 13932 -784 13966
rect -748 13932 -714 13966
rect -678 13932 -644 13966
rect -608 13932 -574 13966
rect -538 13932 -504 13966
rect -468 13932 -434 13966
rect -398 13932 -364 13966
rect -328 13932 -294 13966
rect -258 13932 -224 13966
rect -188 13932 -154 13966
rect -118 13932 -84 13966
rect -48 13932 -14 13966
rect -818 13864 -784 13898
rect -748 13864 -714 13898
rect -678 13864 -644 13898
rect -608 13864 -574 13898
rect -538 13864 -504 13898
rect -468 13864 -434 13898
rect -398 13864 -364 13898
rect -328 13864 -294 13898
rect -258 13864 -224 13898
rect -188 13864 -154 13898
rect -118 13864 -84 13898
rect -48 13864 -14 13898
rect -818 13796 -784 13830
rect -748 13796 -714 13830
rect -678 13796 -644 13830
rect -608 13796 -574 13830
rect -538 13796 -504 13830
rect -468 13796 -434 13830
rect -398 13796 -364 13830
rect -328 13796 -294 13830
rect -258 13796 -224 13830
rect -188 13796 -154 13830
rect -118 13796 -84 13830
rect -48 13796 -14 13830
rect -818 13728 -784 13762
rect -748 13728 -714 13762
rect -678 13728 -644 13762
rect -608 13728 -574 13762
rect -538 13728 -504 13762
rect -468 13728 -434 13762
rect -398 13728 -364 13762
rect -328 13728 -294 13762
rect -258 13728 -224 13762
rect -188 13728 -154 13762
rect -118 13728 -84 13762
rect -48 13728 -14 13762
rect -818 13660 -784 13694
rect -748 13660 -714 13694
rect -678 13660 -644 13694
rect -608 13660 -574 13694
rect -538 13660 -504 13694
rect -468 13660 -434 13694
rect -398 13660 -364 13694
rect -328 13660 -294 13694
rect -258 13660 -224 13694
rect -188 13660 -154 13694
rect -118 13660 -84 13694
rect -48 13660 -14 13694
rect -818 13592 -784 13626
rect -748 13592 -714 13626
rect -678 13592 -644 13626
rect -608 13592 -574 13626
rect -538 13592 -504 13626
rect -468 13592 -434 13626
rect -398 13592 -364 13626
rect -328 13592 -294 13626
rect -258 13592 -224 13626
rect -188 13592 -154 13626
rect -118 13592 -84 13626
rect -48 13592 -14 13626
rect -818 13524 -784 13558
rect -748 13524 -714 13558
rect -678 13524 -644 13558
rect -608 13524 -574 13558
rect -538 13524 -504 13558
rect -468 13524 -434 13558
rect -398 13524 -364 13558
rect -328 13524 -294 13558
rect -258 13524 -224 13558
rect -188 13524 -154 13558
rect -118 13524 -84 13558
rect -48 13524 -14 13558
rect -818 13456 -784 13490
rect -748 13456 -714 13490
rect -678 13456 -644 13490
rect -608 13456 -574 13490
rect -538 13456 -504 13490
rect -468 13456 -434 13490
rect -398 13456 -364 13490
rect -328 13456 -294 13490
rect -258 13456 -224 13490
rect -188 13456 -154 13490
rect -118 13456 -84 13490
rect -48 13456 -14 13490
rect -818 13388 -784 13422
rect -748 13388 -714 13422
rect -678 13388 -644 13422
rect -608 13388 -574 13422
rect -538 13388 -504 13422
rect -468 13388 -434 13422
rect -398 13388 -364 13422
rect -328 13388 -294 13422
rect -258 13388 -224 13422
rect -188 13388 -154 13422
rect -118 13388 -84 13422
rect -48 13388 -14 13422
rect -818 13320 -784 13354
rect -748 13320 -714 13354
rect -678 13320 -644 13354
rect -608 13320 -574 13354
rect -538 13320 -504 13354
rect -468 13320 -434 13354
rect -398 13320 -364 13354
rect -328 13320 -294 13354
rect -258 13320 -224 13354
rect -188 13320 -154 13354
rect -118 13320 -84 13354
rect -48 13320 -14 13354
rect -818 13252 -784 13286
rect -748 13252 -714 13286
rect -678 13252 -644 13286
rect -608 13252 -574 13286
rect -538 13252 -504 13286
rect -468 13252 -434 13286
rect -398 13252 -364 13286
rect -328 13252 -294 13286
rect -258 13252 -224 13286
rect -188 13252 -154 13286
rect -118 13252 -84 13286
rect -48 13252 -14 13286
rect -818 13184 -784 13218
rect -748 13184 -714 13218
rect -678 13184 -644 13218
rect -608 13184 -574 13218
rect -538 13184 -504 13218
rect -468 13184 -434 13218
rect -398 13184 -364 13218
rect -328 13184 -294 13218
rect -258 13184 -224 13218
rect -188 13184 -154 13218
rect -118 13184 -84 13218
rect -48 13184 -14 13218
rect -818 13116 -784 13150
rect -748 13116 -714 13150
rect -678 13116 -644 13150
rect -608 13116 -574 13150
rect -538 13116 -504 13150
rect -468 13116 -434 13150
rect -398 13116 -364 13150
rect -328 13116 -294 13150
rect -258 13116 -224 13150
rect -188 13116 -154 13150
rect -118 13116 -84 13150
rect -48 13116 -14 13150
rect -818 13048 -784 13082
rect -748 13048 -714 13082
rect -678 13048 -644 13082
rect -608 13048 -574 13082
rect -538 13048 -504 13082
rect -468 13048 -434 13082
rect -398 13048 -364 13082
rect -328 13048 -294 13082
rect -258 13048 -224 13082
rect -188 13048 -154 13082
rect -118 13048 -84 13082
rect -48 13048 -14 13082
rect -818 12980 -784 13014
rect -748 12980 -714 13014
rect -678 12980 -644 13014
rect -608 12980 -574 13014
rect -538 12980 -504 13014
rect -468 12980 -434 13014
rect -398 12980 -364 13014
rect -328 12980 -294 13014
rect -258 12980 -224 13014
rect -188 12980 -154 13014
rect -118 12980 -84 13014
rect -48 12980 -14 13014
rect -818 12912 -784 12946
rect -748 12912 -714 12946
rect -678 12912 -644 12946
rect -608 12912 -574 12946
rect -538 12912 -504 12946
rect -468 12912 -434 12946
rect -398 12912 -364 12946
rect -328 12912 -294 12946
rect -258 12912 -224 12946
rect -188 12912 -154 12946
rect -118 12912 -84 12946
rect -48 12912 -14 12946
rect -818 12844 -784 12878
rect -748 12844 -714 12878
rect -678 12844 -644 12878
rect -608 12844 -574 12878
rect -538 12844 -504 12878
rect -468 12844 -434 12878
rect -398 12844 -364 12878
rect -328 12844 -294 12878
rect -258 12844 -224 12878
rect -188 12844 -154 12878
rect -118 12844 -84 12878
rect -48 12844 -14 12878
rect -818 12776 -784 12810
rect -748 12776 -714 12810
rect -678 12776 -644 12810
rect -608 12776 -574 12810
rect -538 12776 -504 12810
rect -468 12776 -434 12810
rect -398 12776 -364 12810
rect -328 12776 -294 12810
rect -258 12776 -224 12810
rect -188 12776 -154 12810
rect -118 12776 -84 12810
rect -48 12776 -14 12810
rect -818 12708 -784 12742
rect -748 12708 -714 12742
rect -678 12708 -644 12742
rect -608 12708 -574 12742
rect -538 12708 -504 12742
rect -468 12708 -434 12742
rect -398 12708 -364 12742
rect -328 12708 -294 12742
rect -258 12708 -224 12742
rect -188 12708 -154 12742
rect -118 12708 -84 12742
rect -48 12708 -14 12742
rect -818 12640 -784 12674
rect -748 12640 -714 12674
rect -678 12640 -644 12674
rect -608 12640 -574 12674
rect -538 12640 -504 12674
rect -468 12640 -434 12674
rect -398 12640 -364 12674
rect -328 12640 -294 12674
rect -258 12640 -224 12674
rect -188 12640 -154 12674
rect -118 12640 -84 12674
rect -48 12640 -14 12674
rect -818 12572 -784 12606
rect -748 12572 -714 12606
rect -678 12572 -644 12606
rect -608 12572 -574 12606
rect -538 12572 -504 12606
rect -468 12572 -434 12606
rect -398 12572 -364 12606
rect -328 12572 -294 12606
rect -258 12572 -224 12606
rect -188 12572 -154 12606
rect -118 12572 -84 12606
rect -48 12572 -14 12606
rect -818 12504 -784 12538
rect -748 12504 -714 12538
rect -678 12504 -644 12538
rect -608 12504 -574 12538
rect -538 12504 -504 12538
rect -468 12504 -434 12538
rect -398 12504 -364 12538
rect -328 12504 -294 12538
rect -258 12504 -224 12538
rect -188 12504 -154 12538
rect -118 12504 -84 12538
rect -48 12504 -14 12538
rect -818 12436 -784 12470
rect -748 12436 -714 12470
rect -678 12436 -644 12470
rect -608 12436 -574 12470
rect -538 12436 -504 12470
rect -468 12436 -434 12470
rect -398 12436 -364 12470
rect -328 12436 -294 12470
rect -258 12436 -224 12470
rect -188 12436 -154 12470
rect -118 12436 -84 12470
rect -48 12436 -14 12470
rect -818 12368 -784 12402
rect -748 12368 -714 12402
rect -678 12368 -644 12402
rect -608 12368 -574 12402
rect -538 12368 -504 12402
rect -468 12368 -434 12402
rect -398 12368 -364 12402
rect -328 12368 -294 12402
rect -258 12368 -224 12402
rect -188 12368 -154 12402
rect -118 12368 -84 12402
rect -48 12368 -14 12402
rect -818 12300 -784 12334
rect -748 12300 -714 12334
rect -678 12300 -644 12334
rect -608 12300 -574 12334
rect -538 12300 -504 12334
rect -468 12300 -434 12334
rect -398 12300 -364 12334
rect -328 12300 -294 12334
rect -258 12300 -224 12334
rect -188 12300 -154 12334
rect -118 12300 -84 12334
rect -48 12300 -14 12334
rect -818 12232 -784 12266
rect -748 12232 -714 12266
rect -678 12232 -644 12266
rect -608 12232 -574 12266
rect -538 12232 -504 12266
rect -468 12232 -434 12266
rect -398 12232 -364 12266
rect -328 12232 -294 12266
rect -258 12232 -224 12266
rect -188 12232 -154 12266
rect -118 12232 -84 12266
rect -48 12232 -14 12266
rect -818 12164 -784 12198
rect -748 12164 -714 12198
rect -678 12164 -644 12198
rect -608 12164 -574 12198
rect -538 12164 -504 12198
rect -468 12164 -434 12198
rect -398 12164 -364 12198
rect -328 12164 -294 12198
rect -258 12164 -224 12198
rect -188 12164 -154 12198
rect -118 12164 -84 12198
rect -48 12164 -14 12198
rect -818 12096 -784 12130
rect -748 12096 -714 12130
rect -678 12096 -644 12130
rect -608 12096 -574 12130
rect -538 12096 -504 12130
rect -468 12096 -434 12130
rect -398 12096 -364 12130
rect -328 12096 -294 12130
rect -258 12096 -224 12130
rect -188 12096 -154 12130
rect -118 12096 -84 12130
rect -48 12096 -14 12130
rect -818 12028 -784 12062
rect -748 12028 -714 12062
rect -678 12028 -644 12062
rect -608 12028 -574 12062
rect -538 12028 -504 12062
rect -468 12028 -434 12062
rect -398 12028 -364 12062
rect -328 12028 -294 12062
rect -258 12028 -224 12062
rect -188 12028 -154 12062
rect -118 12028 -84 12062
rect -48 12028 -14 12062
rect -818 11960 -784 11994
rect -748 11960 -714 11994
rect -678 11960 -644 11994
rect -608 11960 -574 11994
rect -538 11960 -504 11994
rect -468 11960 -434 11994
rect -398 11960 -364 11994
rect -328 11960 -294 11994
rect -258 11960 -224 11994
rect -188 11960 -154 11994
rect -118 11960 -84 11994
rect -48 11960 -14 11994
rect -818 11892 -784 11926
rect -748 11892 -714 11926
rect -678 11892 -644 11926
rect -608 11892 -574 11926
rect -538 11892 -504 11926
rect -468 11892 -434 11926
rect -398 11892 -364 11926
rect -328 11892 -294 11926
rect -258 11892 -224 11926
rect -188 11892 -154 11926
rect -118 11892 -84 11926
rect -48 11892 -14 11926
rect -818 11824 -784 11858
rect -748 11824 -714 11858
rect -678 11824 -644 11858
rect -608 11824 -574 11858
rect -538 11824 -504 11858
rect -468 11824 -434 11858
rect -398 11824 -364 11858
rect -328 11824 -294 11858
rect -258 11824 -224 11858
rect -188 11824 -154 11858
rect -118 11824 -84 11858
rect -48 11824 -14 11858
rect -818 11756 -784 11790
rect -748 11756 -714 11790
rect -678 11756 -644 11790
rect -608 11756 -574 11790
rect -538 11756 -504 11790
rect -468 11756 -434 11790
rect -398 11756 -364 11790
rect -328 11756 -294 11790
rect -258 11756 -224 11790
rect -188 11756 -154 11790
rect -118 11756 -84 11790
rect -48 11756 -14 11790
rect -818 11688 -784 11722
rect -748 11688 -714 11722
rect -678 11688 -644 11722
rect -608 11688 -574 11722
rect -538 11688 -504 11722
rect -468 11688 -434 11722
rect -398 11688 -364 11722
rect -328 11688 -294 11722
rect -258 11688 -224 11722
rect -188 11688 -154 11722
rect -118 11688 -84 11722
rect -48 11688 -14 11722
rect -818 11620 -784 11654
rect -748 11620 -714 11654
rect -678 11620 -644 11654
rect -608 11620 -574 11654
rect -538 11620 -504 11654
rect -468 11620 -434 11654
rect -398 11620 -364 11654
rect -328 11620 -294 11654
rect -258 11620 -224 11654
rect -188 11620 -154 11654
rect -118 11620 -84 11654
rect -48 11620 -14 11654
rect -818 11552 -784 11586
rect -748 11552 -714 11586
rect -678 11552 -644 11586
rect -608 11552 -574 11586
rect -538 11552 -504 11586
rect -468 11552 -434 11586
rect -398 11552 -364 11586
rect -328 11552 -294 11586
rect -258 11552 -224 11586
rect -188 11552 -154 11586
rect -118 11552 -84 11586
rect -48 11552 -14 11586
rect -818 11484 -784 11518
rect -748 11484 -714 11518
rect -678 11484 -644 11518
rect -608 11484 -574 11518
rect -538 11484 -504 11518
rect -468 11484 -434 11518
rect -398 11484 -364 11518
rect -328 11484 -294 11518
rect -258 11484 -224 11518
rect -188 11484 -154 11518
rect -118 11484 -84 11518
rect -48 11484 -14 11518
rect -818 11416 -784 11450
rect -748 11416 -714 11450
rect -678 11416 -644 11450
rect -608 11416 -574 11450
rect -538 11416 -504 11450
rect -468 11416 -434 11450
rect -398 11416 -364 11450
rect -328 11416 -294 11450
rect -258 11416 -224 11450
rect -188 11416 -154 11450
rect -118 11416 -84 11450
rect -48 11416 -14 11450
rect -818 11348 -784 11382
rect -748 11348 -714 11382
rect -678 11348 -644 11382
rect -608 11348 -574 11382
rect -538 11348 -504 11382
rect -468 11348 -434 11382
rect -398 11348 -364 11382
rect -328 11348 -294 11382
rect -258 11348 -224 11382
rect -188 11348 -154 11382
rect -118 11348 -84 11382
rect -48 11348 -14 11382
rect -818 11280 -784 11314
rect -748 11280 -714 11314
rect -678 11280 -644 11314
rect -608 11280 -574 11314
rect -538 11280 -504 11314
rect -468 11280 -434 11314
rect -398 11280 -364 11314
rect -328 11280 -294 11314
rect -258 11280 -224 11314
rect -188 11280 -154 11314
rect -118 11280 -84 11314
rect -48 11280 -14 11314
rect -818 11212 -784 11246
rect -748 11212 -714 11246
rect -678 11212 -644 11246
rect -608 11212 -574 11246
rect -538 11212 -504 11246
rect -468 11212 -434 11246
rect -398 11212 -364 11246
rect -328 11212 -294 11246
rect -258 11212 -224 11246
rect -188 11212 -154 11246
rect -118 11212 -84 11246
rect -48 11212 -14 11246
rect -818 11144 -784 11178
rect -748 11144 -714 11178
rect -678 11144 -644 11178
rect -608 11144 -574 11178
rect -538 11144 -504 11178
rect -468 11144 -434 11178
rect -398 11144 -364 11178
rect -328 11144 -294 11178
rect -258 11144 -224 11178
rect -188 11144 -154 11178
rect -118 11144 -84 11178
rect -48 11144 -14 11178
rect -818 11076 -784 11110
rect -748 11076 -714 11110
rect -678 11076 -644 11110
rect -608 11076 -574 11110
rect -538 11076 -504 11110
rect -468 11076 -434 11110
rect -398 11076 -364 11110
rect -328 11076 -294 11110
rect -258 11076 -224 11110
rect -188 11076 -154 11110
rect -118 11076 -84 11110
rect -48 11076 -14 11110
rect -818 11008 -784 11042
rect -748 11008 -714 11042
rect -678 11008 -644 11042
rect -608 11008 -574 11042
rect -538 11008 -504 11042
rect -468 11008 -434 11042
rect -398 11008 -364 11042
rect -328 11008 -294 11042
rect -258 11008 -224 11042
rect -188 11008 -154 11042
rect -118 11008 -84 11042
rect -48 11008 -14 11042
rect -818 10940 -784 10974
rect -748 10940 -714 10974
rect -678 10940 -644 10974
rect -608 10940 -574 10974
rect -538 10940 -504 10974
rect -468 10940 -434 10974
rect -398 10940 -364 10974
rect -328 10940 -294 10974
rect -258 10940 -224 10974
rect -188 10940 -154 10974
rect -118 10940 -84 10974
rect -48 10940 -14 10974
rect -818 10872 -784 10906
rect -748 10872 -714 10906
rect -678 10872 -644 10906
rect -608 10872 -574 10906
rect -538 10872 -504 10906
rect -468 10872 -434 10906
rect -398 10872 -364 10906
rect -328 10872 -294 10906
rect -258 10872 -224 10906
rect -188 10872 -154 10906
rect -118 10872 -84 10906
rect -48 10872 -14 10906
rect -818 10804 -784 10838
rect -748 10804 -714 10838
rect -678 10804 -644 10838
rect -608 10804 -574 10838
rect -538 10804 -504 10838
rect -468 10804 -434 10838
rect -398 10804 -364 10838
rect -328 10804 -294 10838
rect -258 10804 -224 10838
rect -188 10804 -154 10838
rect -118 10804 -84 10838
rect -48 10804 -14 10838
rect -818 10736 -784 10770
rect -748 10736 -714 10770
rect -678 10736 -644 10770
rect -608 10736 -574 10770
rect -538 10736 -504 10770
rect -468 10736 -434 10770
rect -398 10736 -364 10770
rect -328 10736 -294 10770
rect -258 10736 -224 10770
rect -188 10736 -154 10770
rect -118 10736 -84 10770
rect -48 10736 -14 10770
rect -818 10668 -784 10702
rect -748 10668 -714 10702
rect -678 10668 -644 10702
rect -608 10668 -574 10702
rect -538 10668 -504 10702
rect -468 10668 -434 10702
rect -398 10668 -364 10702
rect -328 10668 -294 10702
rect -258 10668 -224 10702
rect -188 10668 -154 10702
rect -118 10668 -84 10702
rect -48 10668 -14 10702
rect -818 10600 -784 10634
rect -748 10600 -714 10634
rect -678 10600 -644 10634
rect -608 10600 -574 10634
rect -538 10600 -504 10634
rect -468 10600 -434 10634
rect -398 10600 -364 10634
rect -328 10600 -294 10634
rect -258 10600 -224 10634
rect -188 10600 -154 10634
rect -118 10600 -84 10634
rect -48 10600 -14 10634
rect -818 10532 -784 10566
rect -748 10532 -714 10566
rect -678 10532 -644 10566
rect -608 10532 -574 10566
rect -538 10532 -504 10566
rect -468 10532 -434 10566
rect -398 10532 -364 10566
rect -328 10532 -294 10566
rect -258 10532 -224 10566
rect -188 10532 -154 10566
rect -118 10532 -84 10566
rect -48 10532 -14 10566
rect -818 10464 -784 10498
rect -748 10464 -714 10498
rect -678 10464 -644 10498
rect -608 10464 -574 10498
rect -538 10464 -504 10498
rect -468 10464 -434 10498
rect -398 10464 -364 10498
rect -328 10464 -294 10498
rect -258 10464 -224 10498
rect -188 10464 -154 10498
rect -118 10464 -84 10498
rect -48 10464 -14 10498
rect -818 10396 -784 10430
rect -748 10396 -714 10430
rect -678 10396 -644 10430
rect -608 10396 -574 10430
rect -538 10396 -504 10430
rect -468 10396 -434 10430
rect -398 10396 -364 10430
rect -328 10396 -294 10430
rect -258 10396 -224 10430
rect -188 10396 -154 10430
rect -118 10396 -84 10430
rect -48 10396 -14 10430
rect -818 10328 -784 10362
rect -748 10328 -714 10362
rect -678 10328 -644 10362
rect -608 10328 -574 10362
rect -538 10328 -504 10362
rect -468 10328 -434 10362
rect -398 10328 -364 10362
rect -328 10328 -294 10362
rect -258 10328 -224 10362
rect -188 10328 -154 10362
rect -118 10328 -84 10362
rect -48 10328 -14 10362
rect -818 10260 -784 10294
rect -748 10260 -714 10294
rect -678 10260 -644 10294
rect -608 10260 -574 10294
rect -538 10260 -504 10294
rect -468 10260 -434 10294
rect -398 10260 -364 10294
rect -328 10260 -294 10294
rect -258 10260 -224 10294
rect -188 10260 -154 10294
rect -118 10260 -84 10294
rect -48 10260 -14 10294
rect -818 10192 -784 10226
rect -748 10192 -714 10226
rect -678 10192 -644 10226
rect -608 10192 -574 10226
rect -538 10192 -504 10226
rect -468 10192 -434 10226
rect -398 10192 -364 10226
rect -328 10192 -294 10226
rect -258 10192 -224 10226
rect -188 10192 -154 10226
rect -118 10192 -84 10226
rect -48 10192 -14 10226
rect -818 10124 -784 10158
rect -748 10124 -714 10158
rect -678 10124 -644 10158
rect -608 10124 -574 10158
rect -538 10124 -504 10158
rect -468 10124 -434 10158
rect -398 10124 -364 10158
rect -328 10124 -294 10158
rect -258 10124 -224 10158
rect -188 10124 -154 10158
rect -118 10124 -84 10158
rect -48 10124 -14 10158
rect -818 10056 -784 10090
rect -748 10056 -714 10090
rect -678 10056 -644 10090
rect -608 10056 -574 10090
rect -538 10056 -504 10090
rect -468 10056 -434 10090
rect -398 10056 -364 10090
rect -328 10056 -294 10090
rect -258 10056 -224 10090
rect -188 10056 -154 10090
rect -118 10056 -84 10090
rect -48 10056 -14 10090
rect -818 9988 -784 10022
rect -748 9988 -714 10022
rect -678 9988 -644 10022
rect -608 9988 -574 10022
rect -538 9988 -504 10022
rect -468 9988 -434 10022
rect -398 9988 -364 10022
rect -328 9988 -294 10022
rect -258 9988 -224 10022
rect -188 9988 -154 10022
rect -118 9988 -84 10022
rect -48 9988 -14 10022
rect -818 9920 -784 9954
rect -748 9920 -714 9954
rect -678 9920 -644 9954
rect -608 9920 -574 9954
rect -538 9920 -504 9954
rect -468 9920 -434 9954
rect -398 9920 -364 9954
rect -328 9920 -294 9954
rect -258 9920 -224 9954
rect -188 9920 -154 9954
rect -118 9920 -84 9954
rect -48 9920 -14 9954
rect -818 9852 -784 9886
rect -748 9852 -714 9886
rect -678 9852 -644 9886
rect -608 9852 -574 9886
rect -538 9852 -504 9886
rect -468 9852 -434 9886
rect -398 9852 -364 9886
rect -328 9852 -294 9886
rect -258 9852 -224 9886
rect -188 9852 -154 9886
rect -118 9852 -84 9886
rect -48 9852 -14 9886
rect -818 9784 -784 9818
rect -748 9784 -714 9818
rect -678 9784 -644 9818
rect -608 9784 -574 9818
rect -538 9784 -504 9818
rect -468 9784 -434 9818
rect -398 9784 -364 9818
rect -328 9784 -294 9818
rect -258 9784 -224 9818
rect -188 9784 -154 9818
rect -118 9784 -84 9818
rect -48 9784 -14 9818
rect -818 9716 -784 9750
rect -748 9716 -714 9750
rect -678 9716 -644 9750
rect -608 9716 -574 9750
rect -538 9716 -504 9750
rect -468 9716 -434 9750
rect -398 9716 -364 9750
rect -328 9716 -294 9750
rect -258 9716 -224 9750
rect -188 9716 -154 9750
rect -118 9716 -84 9750
rect -48 9716 -14 9750
rect -818 9648 -784 9682
rect -748 9648 -714 9682
rect -678 9648 -644 9682
rect -608 9648 -574 9682
rect -538 9648 -504 9682
rect -468 9648 -434 9682
rect -398 9648 -364 9682
rect -328 9648 -294 9682
rect -258 9648 -224 9682
rect -188 9648 -154 9682
rect -118 9648 -84 9682
rect -48 9648 -14 9682
rect -818 9580 -784 9614
rect -748 9580 -714 9614
rect -678 9580 -644 9614
rect -608 9580 -574 9614
rect -538 9580 -504 9614
rect -468 9580 -434 9614
rect -398 9580 -364 9614
rect -328 9580 -294 9614
rect -258 9580 -224 9614
rect -188 9580 -154 9614
rect -118 9580 -84 9614
rect -48 9580 -14 9614
rect -818 9512 -784 9546
rect -748 9512 -714 9546
rect -678 9512 -644 9546
rect -608 9512 -574 9546
rect -538 9512 -504 9546
rect -468 9512 -434 9546
rect -398 9512 -364 9546
rect -328 9512 -294 9546
rect -258 9512 -224 9546
rect -188 9512 -154 9546
rect -118 9512 -84 9546
rect -48 9512 -14 9546
rect -818 9444 -784 9478
rect -748 9444 -714 9478
rect -678 9444 -644 9478
rect -608 9444 -574 9478
rect -538 9444 -504 9478
rect -468 9444 -434 9478
rect -398 9444 -364 9478
rect -328 9444 -294 9478
rect -258 9444 -224 9478
rect -188 9444 -154 9478
rect -118 9444 -84 9478
rect -48 9444 -14 9478
rect -818 9376 -784 9410
rect -748 9376 -714 9410
rect -678 9376 -644 9410
rect -608 9376 -574 9410
rect -538 9376 -504 9410
rect -468 9376 -434 9410
rect -398 9376 -364 9410
rect -328 9376 -294 9410
rect -258 9376 -224 9410
rect -188 9376 -154 9410
rect -118 9376 -84 9410
rect -48 9376 -14 9410
rect -818 9308 -784 9342
rect -748 9308 -714 9342
rect -678 9308 -644 9342
rect -608 9308 -574 9342
rect -538 9308 -504 9342
rect -468 9308 -434 9342
rect -398 9308 -364 9342
rect -328 9308 -294 9342
rect -258 9308 -224 9342
rect -188 9308 -154 9342
rect -118 9308 -84 9342
rect -48 9308 -14 9342
rect -818 9240 -784 9274
rect -748 9240 -714 9274
rect -678 9240 -644 9274
rect -608 9240 -574 9274
rect -538 9240 -504 9274
rect -468 9240 -434 9274
rect -398 9240 -364 9274
rect -328 9240 -294 9274
rect -258 9240 -224 9274
rect -188 9240 -154 9274
rect -118 9240 -84 9274
rect -48 9240 -14 9274
rect -818 9172 -784 9206
rect -748 9172 -714 9206
rect -678 9172 -644 9206
rect -608 9172 -574 9206
rect -538 9172 -504 9206
rect -468 9172 -434 9206
rect -398 9172 -364 9206
rect -328 9172 -294 9206
rect -258 9172 -224 9206
rect -188 9172 -154 9206
rect -118 9172 -84 9206
rect -48 9172 -14 9206
rect -818 9104 -784 9138
rect -748 9104 -714 9138
rect -678 9104 -644 9138
rect -608 9104 -574 9138
rect -538 9104 -504 9138
rect -468 9104 -434 9138
rect -398 9104 -364 9138
rect -328 9104 -294 9138
rect -258 9104 -224 9138
rect -188 9104 -154 9138
rect -118 9104 -84 9138
rect -48 9104 -14 9138
rect -818 9036 -784 9070
rect -748 9036 -714 9070
rect -678 9036 -644 9070
rect -608 9036 -574 9070
rect -538 9036 -504 9070
rect -468 9036 -434 9070
rect -398 9036 -364 9070
rect -328 9036 -294 9070
rect -258 9036 -224 9070
rect -188 9036 -154 9070
rect -118 9036 -84 9070
rect -48 9036 -14 9070
rect -818 8968 -784 9002
rect -748 8968 -714 9002
rect -678 8968 -644 9002
rect -608 8968 -574 9002
rect -538 8968 -504 9002
rect -468 8968 -434 9002
rect -398 8968 -364 9002
rect -328 8968 -294 9002
rect -258 8968 -224 9002
rect -188 8968 -154 9002
rect -118 8968 -84 9002
rect -48 8968 -14 9002
rect -818 8900 -784 8934
rect -748 8900 -714 8934
rect -678 8900 -644 8934
rect -608 8900 -574 8934
rect -538 8900 -504 8934
rect -468 8900 -434 8934
rect -398 8900 -364 8934
rect -328 8900 -294 8934
rect -258 8900 -224 8934
rect -188 8900 -154 8934
rect -118 8900 -84 8934
rect -48 8900 -14 8934
rect -818 8832 -784 8866
rect -748 8832 -714 8866
rect -678 8832 -644 8866
rect -608 8832 -574 8866
rect -538 8832 -504 8866
rect -468 8832 -434 8866
rect -398 8832 -364 8866
rect -328 8832 -294 8866
rect -258 8832 -224 8866
rect -188 8832 -154 8866
rect -118 8832 -84 8866
rect -48 8832 -14 8866
rect -818 8764 -784 8798
rect -748 8764 -714 8798
rect -678 8764 -644 8798
rect -608 8764 -574 8798
rect -538 8764 -504 8798
rect -468 8764 -434 8798
rect -398 8764 -364 8798
rect -328 8764 -294 8798
rect -258 8764 -224 8798
rect -188 8764 -154 8798
rect -118 8764 -84 8798
rect -48 8764 -14 8798
rect -818 8696 -784 8730
rect -748 8696 -714 8730
rect -678 8696 -644 8730
rect -608 8696 -574 8730
rect -538 8696 -504 8730
rect -468 8696 -434 8730
rect -398 8696 -364 8730
rect -328 8696 -294 8730
rect -258 8696 -224 8730
rect -188 8696 -154 8730
rect -118 8696 -84 8730
rect -48 8696 -14 8730
rect -818 8628 -784 8662
rect -748 8628 -714 8662
rect -678 8628 -644 8662
rect -608 8628 -574 8662
rect -538 8628 -504 8662
rect -468 8628 -434 8662
rect -398 8628 -364 8662
rect -328 8628 -294 8662
rect -258 8628 -224 8662
rect -188 8628 -154 8662
rect -118 8628 -84 8662
rect -48 8628 -14 8662
rect -818 8560 -784 8594
rect -748 8560 -714 8594
rect -678 8560 -644 8594
rect -608 8560 -574 8594
rect -538 8560 -504 8594
rect -468 8560 -434 8594
rect -398 8560 -364 8594
rect -328 8560 -294 8594
rect -258 8560 -224 8594
rect -188 8560 -154 8594
rect -118 8560 -84 8594
rect -48 8560 -14 8594
rect -818 8492 -784 8526
rect -748 8492 -714 8526
rect -678 8492 -644 8526
rect -608 8492 -574 8526
rect -538 8492 -504 8526
rect -468 8492 -434 8526
rect -398 8492 -364 8526
rect -328 8492 -294 8526
rect -258 8492 -224 8526
rect -188 8492 -154 8526
rect -118 8492 -84 8526
rect -48 8492 -14 8526
rect -818 8424 -784 8458
rect -748 8424 -714 8458
rect -678 8424 -644 8458
rect -608 8424 -574 8458
rect -538 8424 -504 8458
rect -468 8424 -434 8458
rect -398 8424 -364 8458
rect -328 8424 -294 8458
rect -258 8424 -224 8458
rect -188 8424 -154 8458
rect -118 8424 -84 8458
rect -48 8424 -14 8458
rect -818 8356 -784 8390
rect -748 8356 -714 8390
rect -678 8356 -644 8390
rect -608 8356 -574 8390
rect -538 8356 -504 8390
rect -468 8356 -434 8390
rect -398 8356 -364 8390
rect -328 8356 -294 8390
rect -258 8356 -224 8390
rect -188 8356 -154 8390
rect -118 8356 -84 8390
rect -48 8356 -14 8390
rect -818 8288 -784 8322
rect -748 8288 -714 8322
rect -678 8288 -644 8322
rect -608 8288 -574 8322
rect -538 8288 -504 8322
rect -468 8288 -434 8322
rect -398 8288 -364 8322
rect -328 8288 -294 8322
rect -258 8288 -224 8322
rect -188 8288 -154 8322
rect -118 8288 -84 8322
rect -48 8288 -14 8322
rect -818 8220 -784 8254
rect -748 8220 -714 8254
rect -678 8220 -644 8254
rect -608 8220 -574 8254
rect -538 8220 -504 8254
rect -468 8220 -434 8254
rect -398 8220 -364 8254
rect -328 8220 -294 8254
rect -258 8220 -224 8254
rect -188 8220 -154 8254
rect -118 8220 -84 8254
rect -48 8220 -14 8254
rect -818 8152 -784 8186
rect -748 8152 -714 8186
rect -678 8152 -644 8186
rect -608 8152 -574 8186
rect -538 8152 -504 8186
rect -468 8152 -434 8186
rect -398 8152 -364 8186
rect -328 8152 -294 8186
rect -258 8152 -224 8186
rect -188 8152 -154 8186
rect -118 8152 -84 8186
rect -48 8152 -14 8186
rect -818 8084 -784 8118
rect -748 8084 -714 8118
rect -678 8084 -644 8118
rect -608 8084 -574 8118
rect -538 8084 -504 8118
rect -468 8084 -434 8118
rect -398 8084 -364 8118
rect -328 8084 -294 8118
rect -258 8084 -224 8118
rect -188 8084 -154 8118
rect -118 8084 -84 8118
rect -48 8084 -14 8118
rect -818 8016 -784 8050
rect -748 8016 -714 8050
rect -678 8016 -644 8050
rect -608 8016 -574 8050
rect -538 8016 -504 8050
rect -468 8016 -434 8050
rect -398 8016 -364 8050
rect -328 8016 -294 8050
rect -258 8016 -224 8050
rect -188 8016 -154 8050
rect -118 8016 -84 8050
rect -48 8016 -14 8050
rect -818 7948 -784 7982
rect -748 7948 -714 7982
rect -678 7948 -644 7982
rect -608 7948 -574 7982
rect -538 7948 -504 7982
rect -468 7948 -434 7982
rect -398 7948 -364 7982
rect -328 7948 -294 7982
rect -258 7948 -224 7982
rect -188 7948 -154 7982
rect -118 7948 -84 7982
rect -48 7948 -14 7982
rect -818 7880 -784 7914
rect -748 7880 -714 7914
rect -678 7880 -644 7914
rect -608 7880 -574 7914
rect -538 7880 -504 7914
rect -468 7880 -434 7914
rect -398 7880 -364 7914
rect -328 7880 -294 7914
rect -258 7880 -224 7914
rect -188 7880 -154 7914
rect -118 7880 -84 7914
rect -48 7880 -14 7914
rect -818 7812 -784 7846
rect -748 7812 -714 7846
rect -678 7812 -644 7846
rect -608 7812 -574 7846
rect -538 7812 -504 7846
rect -468 7812 -434 7846
rect -398 7812 -364 7846
rect -328 7812 -294 7846
rect -258 7812 -224 7846
rect -188 7812 -154 7846
rect -118 7812 -84 7846
rect -48 7812 -14 7846
rect -818 7744 -784 7778
rect -748 7744 -714 7778
rect -678 7744 -644 7778
rect -608 7744 -574 7778
rect -538 7744 -504 7778
rect -468 7744 -434 7778
rect -398 7744 -364 7778
rect -328 7744 -294 7778
rect -258 7744 -224 7778
rect -188 7744 -154 7778
rect -118 7744 -84 7778
rect -48 7744 -14 7778
rect -818 7676 -784 7710
rect -748 7676 -714 7710
rect -678 7676 -644 7710
rect -608 7676 -574 7710
rect -538 7676 -504 7710
rect -468 7676 -434 7710
rect -398 7676 -364 7710
rect -328 7676 -294 7710
rect -258 7676 -224 7710
rect -188 7676 -154 7710
rect -118 7676 -84 7710
rect -48 7676 -14 7710
rect -818 7608 -784 7642
rect -748 7608 -714 7642
rect -678 7608 -644 7642
rect -608 7608 -574 7642
rect -538 7608 -504 7642
rect -468 7608 -434 7642
rect -398 7608 -364 7642
rect -328 7608 -294 7642
rect -258 7608 -224 7642
rect -188 7608 -154 7642
rect -118 7608 -84 7642
rect -48 7608 -14 7642
rect -818 7540 -784 7574
rect -748 7540 -714 7574
rect -678 7540 -644 7574
rect -608 7540 -574 7574
rect -538 7540 -504 7574
rect -468 7540 -434 7574
rect -398 7540 -364 7574
rect -328 7540 -294 7574
rect -258 7540 -224 7574
rect -188 7540 -154 7574
rect -118 7540 -84 7574
rect -48 7540 -14 7574
rect -818 7472 -784 7506
rect -748 7472 -714 7506
rect -678 7472 -644 7506
rect -608 7472 -574 7506
rect -538 7472 -504 7506
rect -468 7472 -434 7506
rect -398 7472 -364 7506
rect -328 7472 -294 7506
rect -258 7472 -224 7506
rect -188 7472 -154 7506
rect -118 7472 -84 7506
rect -48 7472 -14 7506
rect -818 7404 -784 7438
rect -748 7404 -714 7438
rect -678 7404 -644 7438
rect -608 7404 -574 7438
rect -538 7404 -504 7438
rect -468 7404 -434 7438
rect -398 7404 -364 7438
rect -328 7404 -294 7438
rect -258 7404 -224 7438
rect -188 7404 -154 7438
rect -118 7404 -84 7438
rect -48 7404 -14 7438
rect -818 7336 -784 7370
rect -748 7336 -714 7370
rect -678 7336 -644 7370
rect -608 7336 -574 7370
rect -538 7336 -504 7370
rect -468 7336 -434 7370
rect -398 7336 -364 7370
rect -328 7336 -294 7370
rect -258 7336 -224 7370
rect -188 7336 -154 7370
rect -118 7336 -84 7370
rect -48 7336 -14 7370
rect -818 7268 -784 7302
rect -748 7268 -714 7302
rect -678 7268 -644 7302
rect -608 7268 -574 7302
rect -538 7268 -504 7302
rect -468 7268 -434 7302
rect -398 7268 -364 7302
rect -328 7268 -294 7302
rect -258 7268 -224 7302
rect -188 7268 -154 7302
rect -118 7268 -84 7302
rect -48 7268 -14 7302
rect -818 7200 -784 7234
rect -748 7200 -714 7234
rect -678 7200 -644 7234
rect -608 7200 -574 7234
rect -538 7200 -504 7234
rect -468 7200 -434 7234
rect -398 7200 -364 7234
rect -328 7200 -294 7234
rect -258 7200 -224 7234
rect -188 7200 -154 7234
rect -118 7200 -84 7234
rect -48 7200 -14 7234
rect -818 7132 -784 7166
rect -748 7132 -714 7166
rect -678 7132 -644 7166
rect -608 7132 -574 7166
rect -538 7132 -504 7166
rect -468 7132 -434 7166
rect -398 7132 -364 7166
rect -328 7132 -294 7166
rect -258 7132 -224 7166
rect -188 7132 -154 7166
rect -118 7132 -84 7166
rect -48 7132 -14 7166
rect -818 7064 -784 7098
rect -748 7064 -714 7098
rect -678 7064 -644 7098
rect -608 7064 -574 7098
rect -538 7064 -504 7098
rect -468 7064 -434 7098
rect -398 7064 -364 7098
rect -328 7064 -294 7098
rect -258 7064 -224 7098
rect -188 7064 -154 7098
rect -118 7064 -84 7098
rect -48 7064 -14 7098
rect -818 6996 -784 7030
rect -748 6996 -714 7030
rect -678 6996 -644 7030
rect -608 6996 -574 7030
rect -538 6996 -504 7030
rect -468 6996 -434 7030
rect -398 6996 -364 7030
rect -328 6996 -294 7030
rect -258 6996 -224 7030
rect -188 6996 -154 7030
rect -118 6996 -84 7030
rect -48 6996 -14 7030
rect -818 6928 -784 6962
rect -748 6928 -714 6962
rect -678 6928 -644 6962
rect -608 6928 -574 6962
rect -538 6928 -504 6962
rect -468 6928 -434 6962
rect -398 6928 -364 6962
rect -328 6928 -294 6962
rect -258 6928 -224 6962
rect -188 6928 -154 6962
rect -118 6928 -84 6962
rect -48 6928 -14 6962
rect -818 6860 -784 6894
rect -748 6860 -714 6894
rect -678 6860 -644 6894
rect -608 6860 -574 6894
rect -538 6860 -504 6894
rect -468 6860 -434 6894
rect -398 6860 -364 6894
rect -328 6860 -294 6894
rect -258 6860 -224 6894
rect -188 6860 -154 6894
rect -118 6860 -84 6894
rect -48 6860 -14 6894
rect -818 6792 -784 6826
rect -748 6792 -714 6826
rect -678 6792 -644 6826
rect -608 6792 -574 6826
rect -538 6792 -504 6826
rect -468 6792 -434 6826
rect -398 6792 -364 6826
rect -328 6792 -294 6826
rect -258 6792 -224 6826
rect -188 6792 -154 6826
rect -118 6792 -84 6826
rect -48 6792 -14 6826
rect -818 6724 -784 6758
rect -748 6724 -714 6758
rect -678 6724 -644 6758
rect -608 6724 -574 6758
rect -538 6724 -504 6758
rect -468 6724 -434 6758
rect -398 6724 -364 6758
rect -328 6724 -294 6758
rect -258 6724 -224 6758
rect -188 6724 -154 6758
rect -118 6724 -84 6758
rect -48 6724 -14 6758
rect -818 6656 -784 6690
rect -748 6656 -714 6690
rect -678 6656 -644 6690
rect -608 6656 -574 6690
rect -538 6656 -504 6690
rect -468 6656 -434 6690
rect -398 6656 -364 6690
rect -328 6656 -294 6690
rect -258 6656 -224 6690
rect -188 6656 -154 6690
rect -118 6656 -84 6690
rect -48 6656 -14 6690
rect -818 6588 -784 6622
rect -748 6588 -714 6622
rect -678 6588 -644 6622
rect -608 6588 -574 6622
rect -538 6588 -504 6622
rect -468 6588 -434 6622
rect -398 6588 -364 6622
rect -328 6588 -294 6622
rect -258 6588 -224 6622
rect -188 6588 -154 6622
rect -118 6588 -84 6622
rect -48 6588 -14 6622
rect -818 6520 -784 6554
rect -748 6520 -714 6554
rect -678 6520 -644 6554
rect -608 6520 -574 6554
rect -538 6520 -504 6554
rect -468 6520 -434 6554
rect -398 6520 -364 6554
rect -328 6520 -294 6554
rect -258 6520 -224 6554
rect -188 6520 -154 6554
rect -118 6520 -84 6554
rect -48 6520 -14 6554
rect -818 6452 -784 6486
rect -748 6452 -714 6486
rect -678 6452 -644 6486
rect -608 6452 -574 6486
rect -538 6452 -504 6486
rect -468 6452 -434 6486
rect -398 6452 -364 6486
rect -328 6452 -294 6486
rect -258 6452 -224 6486
rect -188 6452 -154 6486
rect -118 6452 -84 6486
rect -48 6452 -14 6486
rect -818 6384 -784 6418
rect -748 6384 -714 6418
rect -678 6384 -644 6418
rect -608 6384 -574 6418
rect -538 6384 -504 6418
rect -468 6384 -434 6418
rect -398 6384 -364 6418
rect -328 6384 -294 6418
rect -258 6384 -224 6418
rect -188 6384 -154 6418
rect -118 6384 -84 6418
rect -48 6384 -14 6418
rect -818 6316 -784 6350
rect -748 6316 -714 6350
rect -678 6316 -644 6350
rect -608 6316 -574 6350
rect -538 6316 -504 6350
rect -468 6316 -434 6350
rect -398 6316 -364 6350
rect -328 6316 -294 6350
rect -258 6316 -224 6350
rect -188 6316 -154 6350
rect -118 6316 -84 6350
rect -48 6316 -14 6350
rect -818 6248 -784 6282
rect -748 6248 -714 6282
rect -678 6248 -644 6282
rect -608 6248 -574 6282
rect -538 6248 -504 6282
rect -468 6248 -434 6282
rect -398 6248 -364 6282
rect -328 6248 -294 6282
rect -258 6248 -224 6282
rect -188 6248 -154 6282
rect -118 6248 -84 6282
rect -48 6248 -14 6282
rect -818 6180 -784 6214
rect -748 6180 -714 6214
rect -678 6180 -644 6214
rect -608 6180 -574 6214
rect -538 6180 -504 6214
rect -468 6180 -434 6214
rect -398 6180 -364 6214
rect -328 6180 -294 6214
rect -258 6180 -224 6214
rect -188 6180 -154 6214
rect -118 6180 -84 6214
rect -48 6180 -14 6214
rect -818 6112 -784 6146
rect -748 6112 -714 6146
rect -678 6112 -644 6146
rect -608 6112 -574 6146
rect -538 6112 -504 6146
rect -468 6112 -434 6146
rect -398 6112 -364 6146
rect -328 6112 -294 6146
rect -258 6112 -224 6146
rect -188 6112 -154 6146
rect -118 6112 -84 6146
rect -48 6112 -14 6146
rect -818 6044 -784 6078
rect -748 6044 -714 6078
rect -678 6044 -644 6078
rect -608 6044 -574 6078
rect -538 6044 -504 6078
rect -468 6044 -434 6078
rect -398 6044 -364 6078
rect -328 6044 -294 6078
rect -258 6044 -224 6078
rect -188 6044 -154 6078
rect -118 6044 -84 6078
rect -48 6044 -14 6078
rect -818 5976 -784 6010
rect -748 5976 -714 6010
rect -678 5976 -644 6010
rect -608 5976 -574 6010
rect -538 5976 -504 6010
rect -468 5976 -434 6010
rect -398 5976 -364 6010
rect -328 5976 -294 6010
rect -258 5976 -224 6010
rect -188 5976 -154 6010
rect -118 5976 -84 6010
rect -48 5976 -14 6010
rect -818 5908 -784 5942
rect -748 5908 -714 5942
rect -678 5908 -644 5942
rect -608 5908 -574 5942
rect -538 5908 -504 5942
rect -468 5908 -434 5942
rect -398 5908 -364 5942
rect -328 5908 -294 5942
rect -258 5908 -224 5942
rect -188 5908 -154 5942
rect -118 5908 -84 5942
rect -48 5908 -14 5942
rect -818 5840 -784 5874
rect -748 5840 -714 5874
rect -678 5840 -644 5874
rect -608 5840 -574 5874
rect -538 5840 -504 5874
rect -468 5840 -434 5874
rect -398 5840 -364 5874
rect -328 5840 -294 5874
rect -258 5840 -224 5874
rect -188 5840 -154 5874
rect -118 5840 -84 5874
rect -48 5840 -14 5874
rect -818 5772 -784 5806
rect -748 5772 -714 5806
rect -678 5772 -644 5806
rect -608 5772 -574 5806
rect -538 5772 -504 5806
rect -468 5772 -434 5806
rect -398 5772 -364 5806
rect -328 5772 -294 5806
rect -258 5772 -224 5806
rect -188 5772 -154 5806
rect -118 5772 -84 5806
rect -48 5772 -14 5806
rect -818 5704 -784 5738
rect -748 5704 -714 5738
rect -678 5704 -644 5738
rect -608 5704 -574 5738
rect -538 5704 -504 5738
rect -468 5704 -434 5738
rect -398 5704 -364 5738
rect -328 5704 -294 5738
rect -258 5704 -224 5738
rect -188 5704 -154 5738
rect -118 5704 -84 5738
rect -48 5704 -14 5738
rect -818 5636 -784 5670
rect -748 5636 -714 5670
rect -678 5636 -644 5670
rect -608 5636 -574 5670
rect -538 5636 -504 5670
rect -468 5636 -434 5670
rect -398 5636 -364 5670
rect -328 5636 -294 5670
rect -258 5636 -224 5670
rect -188 5636 -154 5670
rect -118 5636 -84 5670
rect -48 5636 -14 5670
rect -818 5568 -784 5602
rect -748 5568 -714 5602
rect -678 5568 -644 5602
rect -608 5568 -574 5602
rect -538 5568 -504 5602
rect -468 5568 -434 5602
rect -398 5568 -364 5602
rect -328 5568 -294 5602
rect -258 5568 -224 5602
rect -188 5568 -154 5602
rect -118 5568 -84 5602
rect -48 5568 -14 5602
rect -818 5500 -784 5534
rect -748 5500 -714 5534
rect -678 5500 -644 5534
rect -608 5500 -574 5534
rect -538 5500 -504 5534
rect -468 5500 -434 5534
rect -398 5500 -364 5534
rect -328 5500 -294 5534
rect -258 5500 -224 5534
rect -188 5500 -154 5534
rect -118 5500 -84 5534
rect -48 5500 -14 5534
rect -818 5432 -784 5466
rect -748 5432 -714 5466
rect -678 5432 -644 5466
rect -608 5432 -574 5466
rect -538 5432 -504 5466
rect -468 5432 -434 5466
rect -398 5432 -364 5466
rect -328 5432 -294 5466
rect -258 5432 -224 5466
rect -188 5432 -154 5466
rect -118 5432 -84 5466
rect -48 5432 -14 5466
rect -818 5364 -784 5398
rect -748 5364 -714 5398
rect -678 5364 -644 5398
rect -608 5364 -574 5398
rect -538 5364 -504 5398
rect -468 5364 -434 5398
rect -398 5364 -364 5398
rect -328 5364 -294 5398
rect -258 5364 -224 5398
rect -188 5364 -154 5398
rect -118 5364 -84 5398
rect -48 5364 -14 5398
rect -818 5296 -784 5330
rect -748 5296 -714 5330
rect -678 5296 -644 5330
rect -608 5296 -574 5330
rect -538 5296 -504 5330
rect -468 5296 -434 5330
rect -398 5296 -364 5330
rect -328 5296 -294 5330
rect -258 5296 -224 5330
rect -188 5296 -154 5330
rect -118 5296 -84 5330
rect -48 5296 -14 5330
rect -818 5228 -784 5262
rect -748 5228 -714 5262
rect -678 5228 -644 5262
rect -608 5228 -574 5262
rect -538 5228 -504 5262
rect -468 5228 -434 5262
rect -398 5228 -364 5262
rect -328 5228 -294 5262
rect -258 5228 -224 5262
rect -188 5228 -154 5262
rect -118 5228 -84 5262
rect -48 5228 -14 5262
rect -818 5160 -784 5194
rect -748 5160 -714 5194
rect -678 5160 -644 5194
rect -608 5160 -574 5194
rect -538 5160 -504 5194
rect -468 5160 -434 5194
rect -398 5160 -364 5194
rect -328 5160 -294 5194
rect -258 5160 -224 5194
rect -188 5160 -154 5194
rect -118 5160 -84 5194
rect -48 5160 -14 5194
rect -818 5092 -784 5126
rect -748 5092 -714 5126
rect -678 5092 -644 5126
rect -608 5092 -574 5126
rect -538 5092 -504 5126
rect -468 5092 -434 5126
rect -398 5092 -364 5126
rect -328 5092 -294 5126
rect -258 5092 -224 5126
rect -188 5092 -154 5126
rect -118 5092 -84 5126
rect -48 5092 -14 5126
rect -818 5024 -784 5058
rect -748 5024 -714 5058
rect -678 5024 -644 5058
rect -608 5024 -574 5058
rect -538 5024 -504 5058
rect -468 5024 -434 5058
rect -398 5024 -364 5058
rect -328 5024 -294 5058
rect -258 5024 -224 5058
rect -188 5024 -154 5058
rect -118 5024 -84 5058
rect -48 5024 -14 5058
rect -818 4956 -784 4990
rect -748 4956 -714 4990
rect -678 4956 -644 4990
rect -608 4956 -574 4990
rect -538 4956 -504 4990
rect -468 4956 -434 4990
rect -398 4956 -364 4990
rect -328 4956 -294 4990
rect -258 4956 -224 4990
rect -188 4956 -154 4990
rect -118 4956 -84 4990
rect -48 4956 -14 4990
rect 68 4952 102 4986
rect -818 4888 -784 4922
rect -748 4888 -714 4922
rect -678 4888 -644 4922
rect -608 4888 -574 4922
rect -538 4888 -504 4922
rect -468 4888 -434 4922
rect -398 4888 -364 4922
rect -328 4888 -294 4922
rect -258 4888 -224 4922
rect -188 4888 -154 4922
rect -118 4888 -84 4922
rect -48 4888 -14 4922
rect 68 4884 102 4918
rect -818 4820 -784 4854
rect -748 4820 -714 4854
rect -678 4820 -644 4854
rect -608 4820 -574 4854
rect -538 4820 -504 4854
rect -468 4820 -434 4854
rect -398 4820 -364 4854
rect -328 4820 -294 4854
rect -258 4820 -224 4854
rect -188 4820 -154 4854
rect -118 4820 -84 4854
rect -48 4820 -14 4854
rect 68 4816 102 4850
rect -818 4752 -784 4786
rect -748 4752 -714 4786
rect -678 4752 -644 4786
rect -608 4752 -574 4786
rect -538 4752 -504 4786
rect -468 4752 -434 4786
rect -398 4752 -364 4786
rect -328 4752 -294 4786
rect -258 4752 -224 4786
rect -188 4752 -154 4786
rect -118 4752 -84 4786
rect -48 4752 -14 4786
rect 68 4748 102 4782
rect -818 4684 -784 4718
rect -748 4684 -714 4718
rect -678 4684 -644 4718
rect -608 4684 -574 4718
rect -538 4684 -504 4718
rect -468 4684 -434 4718
rect -398 4684 -364 4718
rect -328 4684 -294 4718
rect -258 4684 -224 4718
rect -188 4684 -154 4718
rect -118 4684 -84 4718
rect -48 4684 -14 4718
rect 68 4680 102 4714
rect -818 4616 -784 4650
rect -748 4616 -714 4650
rect -678 4616 -644 4650
rect -608 4616 -574 4650
rect -538 4616 -504 4650
rect -468 4616 -434 4650
rect -398 4616 -364 4650
rect -328 4616 -294 4650
rect -258 4616 -224 4650
rect -188 4616 -154 4650
rect -118 4616 -84 4650
rect -48 4616 -14 4650
rect 68 4612 102 4646
rect -818 4548 -784 4582
rect -748 4548 -714 4582
rect -678 4548 -644 4582
rect -608 4548 -574 4582
rect -538 4548 -504 4582
rect -468 4548 -434 4582
rect -398 4548 -364 4582
rect -328 4548 -294 4582
rect -258 4548 -224 4582
rect -188 4548 -154 4582
rect -118 4548 -84 4582
rect -48 4548 -14 4582
rect 68 4544 102 4578
rect -818 4480 -784 4514
rect -748 4480 -714 4514
rect -678 4480 -644 4514
rect -608 4480 -574 4514
rect -538 4480 -504 4514
rect -468 4480 -434 4514
rect -398 4480 -364 4514
rect -328 4480 -294 4514
rect -258 4480 -224 4514
rect -188 4480 -154 4514
rect -118 4480 -84 4514
rect -48 4480 -14 4514
rect 68 4476 102 4510
rect -818 4412 -784 4446
rect -748 4412 -714 4446
rect -678 4412 -644 4446
rect -608 4412 -574 4446
rect -538 4412 -504 4446
rect -468 4412 -434 4446
rect -398 4412 -364 4446
rect -328 4412 -294 4446
rect -258 4412 -224 4446
rect -188 4412 -154 4446
rect -118 4412 -84 4446
rect -48 4412 -14 4446
rect 68 4408 102 4442
rect -818 4344 -784 4378
rect -748 4344 -714 4378
rect -678 4344 -644 4378
rect -608 4344 -574 4378
rect -538 4344 -504 4378
rect -468 4344 -434 4378
rect -398 4344 -364 4378
rect -328 4344 -294 4378
rect -258 4344 -224 4378
rect -188 4344 -154 4378
rect -118 4344 -84 4378
rect -48 4344 -14 4378
rect 68 4340 102 4374
rect -818 4276 -784 4310
rect -748 4276 -714 4310
rect -678 4276 -644 4310
rect -608 4276 -574 4310
rect -538 4276 -504 4310
rect -468 4276 -434 4310
rect -398 4276 -364 4310
rect -328 4276 -294 4310
rect -258 4276 -224 4310
rect -188 4276 -154 4310
rect -118 4276 -84 4310
rect -48 4276 -14 4310
rect 68 4272 102 4306
rect -818 4208 -784 4242
rect -748 4208 -714 4242
rect -678 4208 -644 4242
rect -608 4208 -574 4242
rect -538 4208 -504 4242
rect -468 4208 -434 4242
rect -398 4208 -364 4242
rect -328 4208 -294 4242
rect -258 4208 -224 4242
rect -188 4208 -154 4242
rect -118 4208 -84 4242
rect -48 4208 -14 4242
rect 68 4204 102 4238
rect -818 4140 -784 4174
rect -748 4140 -714 4174
rect -678 4140 -644 4174
rect -608 4140 -574 4174
rect -538 4140 -504 4174
rect -468 4140 -434 4174
rect -398 4140 -364 4174
rect -328 4140 -294 4174
rect -258 4140 -224 4174
rect -188 4140 -154 4174
rect -118 4140 -84 4174
rect -48 4140 -14 4174
rect 68 4136 102 4170
rect -818 4072 -784 4106
rect -748 4072 -714 4106
rect -678 4072 -644 4106
rect -608 4072 -574 4106
rect -538 4072 -504 4106
rect -468 4072 -434 4106
rect -398 4072 -364 4106
rect -328 4072 -294 4106
rect -258 4072 -224 4106
rect -188 4072 -154 4106
rect -118 4072 -84 4106
rect -48 4072 -14 4106
rect 68 4068 102 4102
rect -818 4004 -784 4038
rect -748 4004 -714 4038
rect -678 4004 -644 4038
rect -608 4004 -574 4038
rect -538 4004 -504 4038
rect -468 4004 -434 4038
rect -398 4004 -364 4038
rect -328 4004 -294 4038
rect -258 4004 -224 4038
rect -188 4004 -154 4038
rect -118 4004 -84 4038
rect -48 4004 -14 4038
rect 68 4000 102 4034
rect -818 3936 -784 3970
rect -748 3936 -714 3970
rect -678 3936 -644 3970
rect -608 3936 -574 3970
rect -538 3936 -504 3970
rect -468 3936 -434 3970
rect -398 3936 -364 3970
rect -328 3936 -294 3970
rect -258 3936 -224 3970
rect -188 3936 -154 3970
rect -118 3936 -84 3970
rect -48 3936 -14 3970
rect 68 3932 102 3966
rect -818 3868 -784 3902
rect -748 3868 -714 3902
rect -678 3868 -644 3902
rect -608 3868 -574 3902
rect -538 3868 -504 3902
rect -468 3868 -434 3902
rect -398 3868 -364 3902
rect -328 3868 -294 3902
rect -258 3868 -224 3902
rect -188 3868 -154 3902
rect -118 3868 -84 3902
rect -48 3868 -14 3902
rect 68 3864 102 3898
rect -818 3800 -784 3834
rect -748 3800 -714 3834
rect -678 3800 -644 3834
rect -608 3800 -574 3834
rect -538 3800 -504 3834
rect -468 3800 -434 3834
rect -398 3800 -364 3834
rect -328 3800 -294 3834
rect -258 3800 -224 3834
rect -188 3800 -154 3834
rect -118 3800 -84 3834
rect -48 3800 -14 3834
rect 68 3796 102 3830
rect -818 3732 -784 3766
rect -748 3732 -714 3766
rect -678 3732 -644 3766
rect -608 3732 -574 3766
rect -538 3732 -504 3766
rect -468 3732 -434 3766
rect -398 3732 -364 3766
rect -328 3732 -294 3766
rect -258 3732 -224 3766
rect -188 3732 -154 3766
rect -118 3732 -84 3766
rect -48 3732 -14 3766
rect 68 3728 102 3762
rect -818 3664 -784 3698
rect -748 3664 -714 3698
rect -678 3664 -644 3698
rect -608 3664 -574 3698
rect -538 3664 -504 3698
rect -468 3664 -434 3698
rect -398 3664 -364 3698
rect -328 3664 -294 3698
rect -258 3664 -224 3698
rect -188 3664 -154 3698
rect -118 3664 -84 3698
rect -48 3664 -14 3698
rect 68 3660 102 3694
rect -818 3596 -784 3630
rect -748 3596 -714 3630
rect -678 3596 -644 3630
rect -608 3596 -574 3630
rect -538 3596 -504 3630
rect -468 3596 -434 3630
rect -398 3596 -364 3630
rect -328 3596 -294 3630
rect -258 3596 -224 3630
rect -188 3596 -154 3630
rect -118 3596 -84 3630
rect -48 3596 -14 3630
rect 68 3592 102 3626
rect -818 3528 -784 3562
rect -748 3528 -714 3562
rect -678 3528 -644 3562
rect -608 3528 -574 3562
rect -538 3528 -504 3562
rect -468 3528 -434 3562
rect -398 3528 -364 3562
rect -328 3528 -294 3562
rect -258 3528 -224 3562
rect -188 3528 -154 3562
rect -118 3528 -84 3562
rect -48 3528 -14 3562
rect 68 3524 102 3558
rect -818 3460 -784 3494
rect -748 3460 -714 3494
rect -678 3460 -644 3494
rect -608 3460 -574 3494
rect -538 3460 -504 3494
rect -468 3460 -434 3494
rect -398 3460 -364 3494
rect -328 3460 -294 3494
rect -258 3460 -224 3494
rect -188 3460 -154 3494
rect -118 3460 -84 3494
rect -48 3460 -14 3494
rect 68 3456 102 3490
rect -818 3392 -784 3426
rect -748 3392 -714 3426
rect -678 3392 -644 3426
rect -608 3392 -574 3426
rect -538 3392 -504 3426
rect -468 3392 -434 3426
rect -398 3392 -364 3426
rect -328 3392 -294 3426
rect -258 3392 -224 3426
rect -188 3392 -154 3426
rect -118 3392 -84 3426
rect -48 3392 -14 3426
rect 68 3388 102 3422
rect -818 3324 -784 3358
rect -748 3324 -714 3358
rect -678 3324 -644 3358
rect -608 3324 -574 3358
rect -538 3324 -504 3358
rect -468 3324 -434 3358
rect -398 3324 -364 3358
rect -328 3324 -294 3358
rect -258 3324 -224 3358
rect -188 3324 -154 3358
rect -118 3324 -84 3358
rect -48 3324 -14 3358
rect 68 3320 102 3354
rect -818 3256 -784 3290
rect -748 3256 -714 3290
rect -678 3256 -644 3290
rect -608 3256 -574 3290
rect -538 3256 -504 3290
rect -468 3256 -434 3290
rect -398 3256 -364 3290
rect -328 3256 -294 3290
rect -258 3256 -224 3290
rect -188 3256 -154 3290
rect -118 3256 -84 3290
rect -48 3256 -14 3290
rect 68 3252 102 3286
rect -818 3188 -784 3222
rect -748 3188 -714 3222
rect -678 3188 -644 3222
rect -608 3188 -574 3222
rect -538 3188 -504 3222
rect -468 3188 -434 3222
rect -398 3188 -364 3222
rect -328 3188 -294 3222
rect -258 3188 -224 3222
rect -188 3188 -154 3222
rect -118 3188 -84 3222
rect -48 3188 -14 3222
rect 68 3184 102 3218
rect -818 3120 -784 3154
rect -748 3120 -714 3154
rect -678 3120 -644 3154
rect -608 3120 -574 3154
rect -538 3120 -504 3154
rect -468 3120 -434 3154
rect -398 3120 -364 3154
rect -328 3120 -294 3154
rect -258 3120 -224 3154
rect -188 3120 -154 3154
rect -118 3120 -84 3154
rect -48 3120 -14 3154
rect 68 3116 102 3150
rect -818 3052 -784 3086
rect -748 3052 -714 3086
rect -678 3052 -644 3086
rect -608 3052 -574 3086
rect -538 3052 -504 3086
rect -468 3052 -434 3086
rect -398 3052 -364 3086
rect -328 3052 -294 3086
rect -258 3052 -224 3086
rect -188 3052 -154 3086
rect -118 3052 -84 3086
rect -48 3052 -14 3086
rect 68 3048 102 3082
rect -818 2984 -784 3018
rect -748 2984 -714 3018
rect -678 2984 -644 3018
rect -608 2984 -574 3018
rect -538 2984 -504 3018
rect -468 2984 -434 3018
rect -398 2984 -364 3018
rect -328 2984 -294 3018
rect -258 2984 -224 3018
rect -188 2984 -154 3018
rect -118 2984 -84 3018
rect -48 2984 -14 3018
rect 68 2980 102 3014
rect -818 2916 -784 2950
rect -748 2916 -714 2950
rect -678 2916 -644 2950
rect -608 2916 -574 2950
rect -538 2916 -504 2950
rect -468 2916 -434 2950
rect -398 2916 -364 2950
rect -328 2916 -294 2950
rect -258 2916 -224 2950
rect -188 2916 -154 2950
rect -118 2916 -84 2950
rect -48 2916 -14 2950
rect 68 2912 102 2946
rect -818 2848 -784 2882
rect -748 2848 -714 2882
rect -678 2848 -644 2882
rect -608 2848 -574 2882
rect -538 2848 -504 2882
rect -468 2848 -434 2882
rect -398 2848 -364 2882
rect -328 2848 -294 2882
rect -258 2848 -224 2882
rect -188 2848 -154 2882
rect -118 2848 -84 2882
rect -48 2848 -14 2882
rect 68 2844 102 2878
rect -818 2780 -784 2814
rect -748 2780 -714 2814
rect -678 2780 -644 2814
rect -608 2780 -574 2814
rect -538 2780 -504 2814
rect -468 2780 -434 2814
rect -398 2780 -364 2814
rect -328 2780 -294 2814
rect -258 2780 -224 2814
rect -188 2780 -154 2814
rect -118 2780 -84 2814
rect -48 2780 -14 2814
rect 68 2776 102 2810
rect -818 2712 -784 2746
rect -748 2712 -714 2746
rect -678 2712 -644 2746
rect -608 2712 -574 2746
rect -538 2712 -504 2746
rect -468 2712 -434 2746
rect -398 2712 -364 2746
rect -328 2712 -294 2746
rect -258 2712 -224 2746
rect -188 2712 -154 2746
rect -118 2712 -84 2746
rect -48 2712 -14 2746
rect 68 2708 102 2742
rect -818 2644 -784 2678
rect -748 2644 -714 2678
rect -678 2644 -644 2678
rect -608 2644 -574 2678
rect -538 2644 -504 2678
rect -468 2644 -434 2678
rect -398 2644 -364 2678
rect -328 2644 -294 2678
rect -258 2644 -224 2678
rect -188 2644 -154 2678
rect -118 2644 -84 2678
rect -48 2644 -14 2678
rect 68 2640 102 2674
rect -818 2576 -784 2610
rect -748 2576 -714 2610
rect -678 2576 -644 2610
rect -608 2576 -574 2610
rect -538 2576 -504 2610
rect -468 2576 -434 2610
rect -398 2576 -364 2610
rect -328 2576 -294 2610
rect -258 2576 -224 2610
rect -188 2576 -154 2610
rect -118 2576 -84 2610
rect -48 2576 -14 2610
rect 68 2572 102 2606
rect -818 2508 -784 2542
rect -748 2508 -714 2542
rect -678 2508 -644 2542
rect -608 2508 -574 2542
rect -538 2508 -504 2542
rect -468 2508 -434 2542
rect -398 2508 -364 2542
rect -328 2508 -294 2542
rect -258 2508 -224 2542
rect -188 2508 -154 2542
rect -118 2508 -84 2542
rect -48 2508 -14 2542
rect 68 2504 102 2538
rect -818 2439 -784 2473
rect -748 2439 -714 2473
rect -678 2439 -644 2473
rect -608 2439 -574 2473
rect -538 2439 -504 2473
rect -468 2439 -434 2473
rect -398 2439 -364 2473
rect -328 2439 -294 2473
rect -258 2439 -224 2473
rect -188 2439 -154 2473
rect -118 2439 -84 2473
rect -48 2439 -14 2473
rect 68 2436 102 2470
rect -818 2370 -784 2404
rect -748 2370 -714 2404
rect -678 2370 -644 2404
rect -608 2370 -574 2404
rect -538 2370 -504 2404
rect -468 2370 -434 2404
rect -398 2370 -364 2404
rect -328 2370 -294 2404
rect -258 2370 -224 2404
rect -188 2370 -154 2404
rect -118 2370 -84 2404
rect -48 2370 -14 2404
rect 68 2368 102 2402
rect -818 2301 -784 2335
rect -748 2301 -714 2335
rect -678 2301 -644 2335
rect -608 2301 -574 2335
rect -538 2301 -504 2335
rect -468 2301 -434 2335
rect -398 2301 -364 2335
rect -328 2301 -294 2335
rect -258 2301 -224 2335
rect -188 2301 -154 2335
rect -118 2301 -84 2335
rect -48 2301 -14 2335
rect 68 2300 102 2334
rect -818 2232 -784 2266
rect -748 2232 -714 2266
rect -678 2232 -644 2266
rect -608 2232 -574 2266
rect -538 2232 -504 2266
rect -468 2232 -434 2266
rect -398 2232 -364 2266
rect -328 2232 -294 2266
rect -258 2232 -224 2266
rect -188 2232 -154 2266
rect -118 2232 -84 2266
rect -48 2232 -14 2266
rect 68 2232 102 2266
rect -818 2163 -784 2197
rect -748 2163 -714 2197
rect -678 2163 -644 2197
rect -608 2163 -574 2197
rect -538 2163 -504 2197
rect -468 2163 -434 2197
rect -398 2163 -364 2197
rect -328 2163 -294 2197
rect -258 2163 -224 2197
rect -188 2163 -154 2197
rect -118 2163 -84 2197
rect -48 2163 -14 2197
rect 68 2164 102 2198
rect -818 2094 -784 2128
rect -748 2094 -714 2128
rect -678 2094 -644 2128
rect -608 2094 -574 2128
rect -538 2094 -504 2128
rect -468 2094 -434 2128
rect -398 2094 -364 2128
rect -328 2094 -294 2128
rect -258 2094 -224 2128
rect -188 2094 -154 2128
rect -118 2094 -84 2128
rect -48 2094 -14 2128
rect 68 2096 102 2130
rect -818 2025 -784 2059
rect -748 2025 -714 2059
rect -678 2025 -644 2059
rect -608 2025 -574 2059
rect -538 2025 -504 2059
rect -468 2025 -434 2059
rect -398 2025 -364 2059
rect -328 2025 -294 2059
rect -258 2025 -224 2059
rect -188 2025 -154 2059
rect -118 2025 -84 2059
rect -48 2025 -14 2059
rect 68 2028 102 2062
rect -818 1956 -784 1990
rect -748 1956 -714 1990
rect -678 1956 -644 1990
rect -608 1956 -574 1990
rect -538 1956 -504 1990
rect -468 1956 -434 1990
rect -398 1956 -364 1990
rect -328 1956 -294 1990
rect -258 1956 -224 1990
rect -188 1956 -154 1990
rect -118 1956 -84 1990
rect -48 1956 -14 1990
rect 68 1960 102 1994
rect -818 1887 -784 1921
rect -748 1887 -714 1921
rect -678 1887 -644 1921
rect -608 1887 -574 1921
rect -538 1887 -504 1921
rect -468 1887 -434 1921
rect -398 1887 -364 1921
rect -328 1887 -294 1921
rect -258 1887 -224 1921
rect -188 1887 -154 1921
rect -118 1887 -84 1921
rect -48 1887 -14 1921
rect 68 1892 102 1926
rect -818 1818 -784 1852
rect -748 1818 -714 1852
rect -678 1818 -644 1852
rect -608 1818 -574 1852
rect -538 1818 -504 1852
rect -468 1818 -434 1852
rect -398 1818 -364 1852
rect -328 1818 -294 1852
rect -258 1818 -224 1852
rect -188 1818 -154 1852
rect -118 1818 -84 1852
rect -48 1818 -14 1852
rect 68 1824 102 1858
rect -818 1749 -784 1783
rect -748 1749 -714 1783
rect -678 1749 -644 1783
rect -608 1749 -574 1783
rect -538 1749 -504 1783
rect -468 1749 -434 1783
rect -398 1749 -364 1783
rect -328 1749 -294 1783
rect -258 1749 -224 1783
rect -188 1749 -154 1783
rect -118 1749 -84 1783
rect -48 1749 -14 1783
rect 68 1756 102 1790
rect -818 1680 -784 1714
rect -748 1680 -714 1714
rect -678 1680 -644 1714
rect -608 1680 -574 1714
rect -538 1680 -504 1714
rect -468 1680 -434 1714
rect -398 1680 -364 1714
rect -328 1680 -294 1714
rect -258 1680 -224 1714
rect -188 1680 -154 1714
rect -118 1680 -84 1714
rect -48 1680 -14 1714
rect 68 1688 102 1722
rect -818 1611 -784 1645
rect -748 1611 -714 1645
rect -678 1611 -644 1645
rect -608 1611 -574 1645
rect -538 1611 -504 1645
rect -468 1611 -434 1645
rect -398 1611 -364 1645
rect -328 1611 -294 1645
rect -258 1611 -224 1645
rect -188 1611 -154 1645
rect -118 1611 -84 1645
rect -48 1611 -14 1645
rect 68 1620 102 1654
rect -818 1542 -784 1576
rect -748 1542 -714 1576
rect -678 1542 -644 1576
rect -608 1542 -574 1576
rect -538 1542 -504 1576
rect -468 1542 -434 1576
rect -398 1542 -364 1576
rect -328 1542 -294 1576
rect -258 1542 -224 1576
rect -188 1542 -154 1576
rect -118 1542 -84 1576
rect -48 1542 -14 1576
rect 68 1552 102 1586
rect -818 1473 -784 1507
rect -748 1473 -714 1507
rect -678 1473 -644 1507
rect -608 1473 -574 1507
rect -538 1473 -504 1507
rect -468 1473 -434 1507
rect -398 1473 -364 1507
rect -328 1473 -294 1507
rect -258 1473 -224 1507
rect -188 1473 -154 1507
rect -118 1473 -84 1507
rect -48 1473 -14 1507
rect 68 1484 102 1518
rect -818 1404 -784 1438
rect -748 1404 -714 1438
rect -678 1404 -644 1438
rect -608 1404 -574 1438
rect -538 1404 -504 1438
rect -468 1404 -434 1438
rect -398 1404 -364 1438
rect -328 1404 -294 1438
rect -258 1404 -224 1438
rect -188 1404 -154 1438
rect -118 1404 -84 1438
rect -48 1404 -14 1438
rect 68 1416 102 1450
rect -818 1335 -784 1369
rect -748 1335 -714 1369
rect -678 1335 -644 1369
rect -608 1335 -574 1369
rect -538 1335 -504 1369
rect -468 1335 -434 1369
rect -398 1335 -364 1369
rect -328 1335 -294 1369
rect -258 1335 -224 1369
rect -188 1335 -154 1369
rect -118 1335 -84 1369
rect -48 1335 -14 1369
rect 68 1347 102 1381
rect -818 1266 -784 1300
rect -748 1266 -714 1300
rect -678 1266 -644 1300
rect -608 1266 -574 1300
rect -538 1266 -504 1300
rect -468 1266 -434 1300
rect -398 1266 -364 1300
rect -328 1266 -294 1300
rect -258 1266 -224 1300
rect -188 1266 -154 1300
rect -118 1266 -84 1300
rect -48 1266 -14 1300
rect 68 1278 102 1312
rect -818 1197 -784 1231
rect -748 1197 -714 1231
rect -678 1197 -644 1231
rect -608 1197 -574 1231
rect -538 1197 -504 1231
rect -468 1197 -434 1231
rect -398 1197 -364 1231
rect -328 1197 -294 1231
rect -258 1197 -224 1231
rect -188 1197 -154 1231
rect -118 1197 -84 1231
rect -48 1197 -14 1231
rect 68 1209 102 1243
rect -818 1128 -784 1162
rect -748 1128 -714 1162
rect -678 1128 -644 1162
rect -608 1128 -574 1162
rect -538 1128 -504 1162
rect -468 1128 -434 1162
rect -398 1128 -364 1162
rect -328 1128 -294 1162
rect -258 1128 -224 1162
rect -188 1128 -154 1162
rect -118 1128 -84 1162
rect -48 1128 -14 1162
rect 68 1140 102 1174
rect -818 1059 -784 1093
rect -748 1059 -714 1093
rect -678 1059 -644 1093
rect -608 1059 -574 1093
rect -538 1059 -504 1093
rect -468 1059 -434 1093
rect -398 1059 -364 1093
rect -328 1059 -294 1093
rect -258 1059 -224 1093
rect -188 1059 -154 1093
rect -118 1059 -84 1093
rect -48 1059 -14 1093
rect 68 1071 102 1105
rect -818 990 -784 1024
rect -748 990 -714 1024
rect -678 990 -644 1024
rect -608 990 -574 1024
rect -538 990 -504 1024
rect -468 990 -434 1024
rect -398 990 -364 1024
rect -328 990 -294 1024
rect -258 990 -224 1024
rect -188 990 -154 1024
rect -118 990 -84 1024
rect -48 990 -14 1024
rect 68 1002 102 1036
rect -818 921 -784 955
rect -748 921 -714 955
rect -678 921 -644 955
rect -608 921 -574 955
rect -538 921 -504 955
rect -468 921 -434 955
rect -398 921 -364 955
rect -328 921 -294 955
rect -258 921 -224 955
rect -188 921 -154 955
rect -118 921 -84 955
rect -48 921 -14 955
rect 68 933 102 967
rect -818 852 -784 886
rect -748 852 -714 886
rect -678 852 -644 886
rect -608 852 -574 886
rect -538 852 -504 886
rect -468 852 -434 886
rect -398 852 -364 886
rect -328 852 -294 886
rect -258 852 -224 886
rect -188 852 -154 886
rect -118 852 -84 886
rect -48 852 -14 886
rect 68 864 102 898
rect -818 783 -784 817
rect -748 783 -714 817
rect -678 783 -644 817
rect -608 783 -574 817
rect -538 783 -504 817
rect -468 783 -434 817
rect -398 783 -364 817
rect -328 783 -294 817
rect -258 783 -224 817
rect -188 783 -154 817
rect -118 783 -84 817
rect -48 783 -14 817
rect 68 795 102 829
rect -818 714 -784 748
rect -748 714 -714 748
rect -678 714 -644 748
rect -608 714 -574 748
rect -538 714 -504 748
rect -468 714 -434 748
rect -398 714 -364 748
rect -328 714 -294 748
rect -258 714 -224 748
rect -188 714 -154 748
rect -118 714 -84 748
rect -48 714 -14 748
rect 68 726 102 760
rect -818 645 -784 679
rect -748 645 -714 679
rect -678 645 -644 679
rect -608 645 -574 679
rect -538 645 -504 679
rect -468 645 -434 679
rect -398 645 -364 679
rect -328 645 -294 679
rect -258 645 -224 679
rect -188 645 -154 679
rect -118 645 -84 679
rect -48 645 -14 679
rect 68 657 102 691
rect -818 576 -784 610
rect -748 576 -714 610
rect -678 576 -644 610
rect -608 576 -574 610
rect -538 576 -504 610
rect -468 576 -434 610
rect -398 576 -364 610
rect -328 576 -294 610
rect -258 576 -224 610
rect -188 576 -154 610
rect -118 576 -84 610
rect -48 576 -14 610
rect 68 588 102 622
rect -818 507 -784 541
rect -748 507 -714 541
rect -678 507 -644 541
rect -608 507 -574 541
rect -538 507 -504 541
rect -468 507 -434 541
rect -398 507 -364 541
rect -328 507 -294 541
rect -258 507 -224 541
rect -188 507 -154 541
rect -118 507 -84 541
rect -48 507 -14 541
rect 68 519 102 553
rect -818 438 -784 472
rect -748 438 -714 472
rect -678 438 -644 472
rect -608 438 -574 472
rect -538 438 -504 472
rect -468 438 -434 472
rect -398 438 -364 472
rect -328 438 -294 472
rect -258 438 -224 472
rect -188 438 -154 472
rect -118 438 -84 472
rect -48 438 -14 472
rect 68 450 102 484
rect -818 369 -784 403
rect -748 369 -714 403
rect -678 369 -644 403
rect -608 369 -574 403
rect -538 369 -504 403
rect -468 369 -434 403
rect -398 369 -364 403
rect -328 369 -294 403
rect -258 369 -224 403
rect -188 369 -154 403
rect -118 369 -84 403
rect -48 369 -14 403
rect 68 381 102 415
rect -818 300 -784 334
rect -748 300 -714 334
rect -678 300 -644 334
rect -608 300 -574 334
rect -538 300 -504 334
rect -468 300 -434 334
rect -398 300 -364 334
rect -328 300 -294 334
rect -258 300 -224 334
rect -188 300 -154 334
rect -118 300 -84 334
rect -48 300 -14 334
rect 68 312 102 346
rect -818 231 -784 265
rect -748 231 -714 265
rect -678 231 -644 265
rect -608 231 -574 265
rect -538 231 -504 265
rect -468 231 -434 265
rect -398 231 -364 265
rect -328 231 -294 265
rect -258 231 -224 265
rect -188 231 -154 265
rect -118 231 -84 265
rect -48 231 -14 265
rect 68 243 102 277
rect -818 162 -784 196
rect -748 162 -714 196
rect -678 162 -644 196
rect -608 162 -574 196
rect -538 162 -504 196
rect -468 162 -434 196
rect -398 162 -364 196
rect -328 162 -294 196
rect -258 162 -224 196
rect -188 162 -154 196
rect -118 162 -84 196
rect -48 162 -14 196
rect 68 174 102 208
rect -818 93 -784 127
rect -748 93 -714 127
rect -678 93 -644 127
rect -608 93 -574 127
rect -538 93 -504 127
rect -468 93 -434 127
rect -398 93 -364 127
rect -328 93 -294 127
rect -258 93 -224 127
rect -188 93 -154 127
rect -118 93 -84 127
rect -48 93 -14 127
rect 92 68 126 102
rect 161 68 195 102
rect 230 68 264 102
rect 300 68 334 102
rect 370 68 404 102
rect 440 68 474 102
rect 510 68 544 102
rect 580 68 614 102
rect 650 68 684 102
rect 720 68 754 102
rect 790 68 824 102
rect -818 24 -784 58
rect -748 24 -714 58
rect -678 24 -644 58
rect -608 24 -574 58
rect -538 24 -504 58
rect -468 24 -434 58
rect -398 24 -364 58
rect -328 24 -294 58
rect -258 24 -224 58
rect -188 24 -154 58
rect -118 24 -84 58
rect -48 24 -14 58
rect 92 0 126 34
rect 161 0 195 34
rect 230 0 264 34
rect 300 0 334 34
rect 370 0 404 34
rect 440 0 474 34
rect 510 0 544 34
rect 580 0 614 34
rect 650 0 684 34
rect 720 0 754 34
rect 790 0 824 34
rect -818 -68 -784 -34
rect -750 -68 -716 -34
rect -682 -68 -648 -34
rect -614 -68 -580 -34
rect -546 -68 -512 -34
rect -478 -68 -444 -34
rect -410 -68 -376 -34
rect -342 -68 -308 -34
rect -274 -68 -240 -34
rect -205 -68 -171 -34
rect -136 -68 -102 -34
rect -67 -68 -33 -34
rect 2 -68 36 -34
rect 71 -68 105 -34
rect 140 -68 174 -34
rect 209 -68 243 -34
rect 278 -68 312 -34
rect 347 -68 381 -34
rect 416 -68 450 -34
rect 485 -68 519 -34
rect 554 -68 588 -34
rect 623 -68 657 -34
rect 692 -68 726 -34
rect 761 -68 795 -34
rect 830 -68 864 -34
rect -818 -139 -784 -105
rect -750 -139 -716 -105
rect -682 -139 -648 -105
rect -614 -139 -580 -105
rect -546 -139 -512 -105
rect -478 -139 -444 -105
rect -410 -139 -376 -105
rect -342 -139 -308 -105
rect -274 -139 -240 -105
rect -205 -139 -171 -105
rect -136 -139 -102 -105
rect -67 -139 -33 -105
rect 2 -139 36 -105
rect 71 -139 105 -105
rect 140 -139 174 -105
rect 209 -139 243 -105
rect 278 -139 312 -105
rect 347 -139 381 -105
rect 416 -139 450 -105
rect 485 -139 519 -105
rect 554 -139 588 -105
rect 623 -139 657 -105
rect 692 -139 726 -105
rect 761 -139 795 -105
rect 830 -139 864 -105
rect -818 -210 -784 -176
rect -750 -210 -716 -176
rect -682 -210 -648 -176
rect -614 -210 -580 -176
rect -546 -210 -512 -176
rect -478 -210 -444 -176
rect -410 -210 -376 -176
rect -342 -210 -308 -176
rect -274 -210 -240 -176
rect -205 -210 -171 -176
rect -136 -210 -102 -176
rect -67 -210 -33 -176
rect 2 -210 36 -176
rect 71 -210 105 -176
rect 140 -210 174 -176
rect 209 -210 243 -176
rect 278 -210 312 -176
rect 347 -210 381 -176
rect 416 -210 450 -176
rect 485 -210 519 -176
rect 554 -210 588 -176
rect 623 -210 657 -176
rect 692 -210 726 -176
rect 761 -210 795 -176
rect 830 -210 864 -176
rect -818 -281 -784 -247
rect -750 -281 -716 -247
rect -682 -281 -648 -247
rect -614 -281 -580 -247
rect -546 -281 -512 -247
rect -478 -281 -444 -247
rect -410 -281 -376 -247
rect -342 -281 -308 -247
rect -274 -281 -240 -247
rect -205 -281 -171 -247
rect -136 -281 -102 -247
rect -67 -281 -33 -247
rect 2 -281 36 -247
rect 71 -281 105 -247
rect 140 -281 174 -247
rect 209 -281 243 -247
rect 278 -281 312 -247
rect 347 -281 381 -247
rect 416 -281 450 -247
rect 485 -281 519 -247
rect 554 -281 588 -247
rect 623 -281 657 -247
rect 692 -281 726 -247
rect 761 -281 795 -247
rect 830 -281 864 -247
rect -818 -352 -784 -318
rect -750 -352 -716 -318
rect -682 -352 -648 -318
rect -614 -352 -580 -318
rect -546 -352 -512 -318
rect -478 -352 -444 -318
rect -410 -352 -376 -318
rect -342 -352 -308 -318
rect -274 -352 -240 -318
rect -205 -352 -171 -318
rect -136 -352 -102 -318
rect -67 -352 -33 -318
rect 2 -352 36 -318
rect 71 -352 105 -318
rect 140 -352 174 -318
rect 209 -352 243 -318
rect 278 -352 312 -318
rect 347 -352 381 -318
rect 416 -352 450 -318
rect 485 -352 519 -318
rect 554 -352 588 -318
rect 623 -352 657 -318
rect 692 -352 726 -318
rect 761 -352 795 -318
rect 830 -352 864 -318
<< poly >>
rect 415 4714 535 4740
rect 415 3674 535 3714
rect 415 3640 472 3674
rect 506 3640 535 3674
rect 415 3593 535 3640
rect 415 2553 535 2593
rect 415 2519 472 2553
rect 506 2519 535 2553
rect 415 2472 535 2519
rect 415 1434 535 1472
rect 415 1400 472 1434
rect 506 1400 535 1434
rect 415 1362 535 1400
rect 415 336 535 362
<< polycont >>
rect 472 3640 506 3674
rect 472 2519 506 2553
rect 472 1400 506 1434
<< locali >>
rect -852 14682 898 14686
rect -852 14648 -828 14682
rect -794 14648 -759 14682
rect -725 14648 -690 14682
rect -656 14648 -621 14682
rect -587 14648 -552 14682
rect -518 14648 -483 14682
rect -449 14648 -414 14682
rect -380 14648 -345 14682
rect -311 14648 -276 14682
rect -242 14648 -207 14682
rect -173 14648 -138 14682
rect -104 14648 -69 14682
rect -35 14648 0 14682
rect 34 14648 69 14682
rect 103 14648 138 14682
rect 172 14648 207 14682
rect 241 14648 276 14682
rect 310 14648 345 14682
rect 379 14648 414 14682
rect 448 14648 483 14682
rect 517 14648 552 14682
rect 586 14648 621 14682
rect 655 14648 690 14682
rect 724 14648 759 14682
rect 793 14648 828 14682
rect 862 14648 898 14682
rect -852 14610 898 14648
rect -852 14576 -828 14610
rect -794 14576 -759 14610
rect -725 14576 -690 14610
rect -656 14576 -621 14610
rect -587 14576 -552 14610
rect -518 14576 -483 14610
rect -449 14576 -414 14610
rect -380 14576 -345 14610
rect -311 14576 -276 14610
rect -242 14576 -207 14610
rect -173 14576 -138 14610
rect -104 14576 -69 14610
rect -35 14576 0 14610
rect 34 14576 69 14610
rect 103 14576 138 14610
rect 172 14576 207 14610
rect 241 14576 276 14610
rect 310 14576 345 14610
rect 379 14576 414 14610
rect 448 14576 483 14610
rect 517 14576 552 14610
rect 586 14576 621 14610
rect 655 14576 690 14610
rect 724 14576 759 14610
rect 793 14576 828 14610
rect 862 14576 898 14610
rect -852 14538 898 14576
rect -852 14504 -828 14538
rect -794 14517 -759 14538
rect -784 14504 -759 14517
rect -725 14504 -690 14538
rect -656 14504 -621 14538
rect -587 14504 -552 14538
rect -518 14504 -483 14538
rect -449 14504 -414 14538
rect -380 14504 -345 14538
rect -311 14505 -276 14538
rect -242 14505 -207 14538
rect -173 14505 -138 14538
rect -311 14504 -305 14505
rect -242 14504 -231 14505
rect -173 14504 -157 14505
rect -104 14504 -69 14538
rect -35 14504 0 14538
rect 34 14504 69 14538
rect 103 14504 138 14538
rect 172 14504 207 14538
rect 241 14504 276 14538
rect 310 14504 345 14538
rect 379 14504 414 14538
rect 448 14504 483 14538
rect 517 14504 552 14538
rect 586 14504 621 14538
rect 655 14504 690 14538
rect 724 14504 759 14538
rect 793 14504 828 14538
rect 862 14504 898 14538
rect -852 14483 -818 14504
rect -784 14483 -305 14504
rect -852 14471 -305 14483
rect -271 14471 -231 14504
rect -197 14471 -157 14504
rect -123 14471 898 14504
rect -852 14466 898 14471
rect -852 14432 -828 14466
rect -794 14445 -759 14466
rect -784 14432 -759 14445
rect -725 14432 -690 14466
rect -656 14432 -621 14466
rect -587 14432 -552 14466
rect -518 14432 -483 14466
rect -449 14432 -414 14466
rect -380 14432 -345 14466
rect -311 14433 -276 14466
rect -242 14433 -207 14466
rect -173 14433 -138 14466
rect -311 14432 -305 14433
rect -242 14432 -231 14433
rect -173 14432 -157 14433
rect -104 14432 -69 14466
rect -35 14432 0 14466
rect 34 14432 69 14466
rect 103 14432 138 14466
rect 172 14432 207 14466
rect 241 14462 276 14466
rect 310 14462 345 14466
rect 379 14462 414 14466
rect 245 14432 276 14462
rect 327 14432 345 14462
rect 409 14432 414 14462
rect 448 14462 483 14466
rect 517 14462 552 14466
rect 448 14432 457 14462
rect 517 14432 539 14462
rect 586 14432 621 14466
rect 655 14432 690 14466
rect 724 14462 759 14466
rect 737 14432 759 14462
rect 793 14432 828 14466
rect 862 14432 898 14466
rect -852 14411 -818 14432
rect -784 14411 -305 14432
rect -852 14399 -305 14411
rect -271 14399 -231 14432
rect -197 14399 -157 14432
rect -123 14428 211 14432
rect 245 14428 293 14432
rect 327 14428 375 14432
rect 409 14428 457 14432
rect 491 14428 539 14432
rect 573 14428 621 14432
rect 655 14428 703 14432
rect 737 14428 898 14432
rect -123 14399 898 14428
rect -852 14394 898 14399
rect -852 14360 -828 14394
rect -794 14373 -759 14394
rect -784 14360 -759 14373
rect -725 14360 -690 14394
rect -656 14360 -621 14394
rect -587 14360 -552 14394
rect -518 14360 -483 14394
rect -449 14360 -414 14394
rect -380 14360 -345 14394
rect -311 14361 -276 14394
rect -242 14361 -207 14394
rect -173 14361 -138 14394
rect -311 14360 -305 14361
rect -242 14360 -231 14361
rect -173 14360 -157 14361
rect -104 14360 -69 14394
rect -35 14360 0 14394
rect 34 14360 69 14394
rect 103 14360 138 14394
rect 172 14360 207 14394
rect 241 14389 276 14394
rect 310 14389 345 14394
rect 379 14389 414 14394
rect 245 14360 276 14389
rect 327 14360 345 14389
rect 409 14360 414 14389
rect 448 14389 483 14394
rect 517 14389 552 14394
rect 448 14360 457 14389
rect 517 14360 539 14389
rect 586 14360 621 14394
rect 655 14360 690 14394
rect 724 14389 759 14394
rect 737 14360 759 14389
rect 793 14360 828 14394
rect 862 14360 898 14394
rect -852 14339 -818 14360
rect -784 14339 -305 14360
rect -852 14327 -305 14339
rect -271 14327 -231 14360
rect -197 14327 -157 14360
rect -123 14355 211 14360
rect 245 14355 293 14360
rect 327 14355 375 14360
rect 409 14355 457 14360
rect 491 14355 539 14360
rect 573 14355 621 14360
rect 655 14355 703 14360
rect 737 14355 898 14360
rect -123 14327 898 14355
rect -852 14322 898 14327
rect -852 14288 -828 14322
rect -794 14301 -759 14322
rect -784 14288 -759 14301
rect -725 14288 -690 14322
rect -656 14288 -621 14322
rect -587 14288 -552 14322
rect -518 14288 -483 14322
rect -449 14288 -414 14322
rect -380 14288 -345 14322
rect -311 14289 -276 14322
rect -242 14289 -207 14322
rect -173 14289 -138 14322
rect -311 14288 -305 14289
rect -242 14288 -231 14289
rect -173 14288 -157 14289
rect -104 14288 -69 14322
rect -35 14288 0 14322
rect 34 14288 69 14322
rect 103 14288 138 14322
rect 172 14288 207 14322
rect 241 14316 276 14322
rect 310 14316 345 14322
rect 379 14316 414 14322
rect 245 14288 276 14316
rect 327 14288 345 14316
rect 409 14288 414 14316
rect 448 14316 483 14322
rect 517 14316 552 14322
rect 448 14288 457 14316
rect 517 14288 539 14316
rect 586 14288 621 14322
rect 655 14288 690 14322
rect 724 14316 759 14322
rect 737 14288 759 14316
rect 793 14288 828 14322
rect 862 14288 898 14322
rect -852 14267 -818 14288
rect -784 14267 -305 14288
rect -852 14255 -305 14267
rect -271 14255 -231 14288
rect -197 14255 -157 14288
rect -123 14282 211 14288
rect 245 14282 293 14288
rect 327 14282 375 14288
rect 409 14282 457 14288
rect 491 14282 539 14288
rect 573 14282 621 14288
rect 655 14282 703 14288
rect 737 14282 898 14288
rect -123 14255 898 14282
rect -852 14250 898 14255
rect -852 14216 -828 14250
rect -794 14229 -759 14250
rect -784 14216 -759 14229
rect -725 14216 -690 14250
rect -656 14216 -621 14250
rect -587 14216 -552 14250
rect -518 14216 -483 14250
rect -449 14216 -414 14250
rect -380 14216 -345 14250
rect -311 14217 -276 14250
rect -242 14217 -207 14250
rect -173 14217 -138 14250
rect -311 14216 -305 14217
rect -242 14216 -231 14217
rect -173 14216 -157 14217
rect -104 14216 -69 14250
rect -35 14216 0 14250
rect 34 14216 69 14250
rect 103 14216 138 14250
rect 172 14216 207 14250
rect 241 14243 276 14250
rect 310 14243 345 14250
rect 379 14243 414 14250
rect 245 14216 276 14243
rect 327 14216 345 14243
rect 409 14216 414 14243
rect 448 14243 483 14250
rect 517 14243 552 14250
rect 448 14216 457 14243
rect 517 14216 539 14243
rect 586 14216 621 14250
rect 655 14216 690 14250
rect 724 14243 759 14250
rect 737 14216 759 14243
rect 793 14216 828 14250
rect 862 14216 898 14250
rect -852 14195 -818 14216
rect -784 14195 -305 14216
rect -852 14183 -305 14195
rect -271 14183 -231 14216
rect -197 14183 -157 14216
rect -123 14209 211 14216
rect 245 14209 293 14216
rect 327 14209 375 14216
rect 409 14209 457 14216
rect 491 14209 539 14216
rect 573 14209 621 14216
rect 655 14209 703 14216
rect 737 14209 898 14216
rect -123 14183 898 14209
rect -852 14178 898 14183
rect -852 14144 -828 14178
rect -794 14157 -759 14178
rect -784 14144 -759 14157
rect -725 14144 -690 14178
rect -656 14144 -621 14178
rect -587 14144 -552 14178
rect -518 14144 -483 14178
rect -449 14144 -414 14178
rect -380 14144 -345 14178
rect -311 14145 -276 14178
rect -242 14145 -207 14178
rect -173 14145 -138 14178
rect -311 14144 -305 14145
rect -242 14144 -231 14145
rect -173 14144 -157 14145
rect -104 14144 -69 14178
rect -35 14144 0 14178
rect 34 14144 69 14178
rect 103 14144 138 14178
rect 172 14144 207 14178
rect 241 14170 276 14178
rect 310 14170 345 14178
rect 379 14170 414 14178
rect 245 14144 276 14170
rect 327 14144 345 14170
rect 409 14144 414 14170
rect 448 14170 483 14178
rect 517 14170 552 14178
rect 448 14144 457 14170
rect 517 14144 539 14170
rect 586 14144 621 14178
rect 655 14144 690 14178
rect 724 14170 759 14178
rect 737 14144 759 14170
rect 793 14144 828 14178
rect 862 14144 898 14178
rect -852 14123 -818 14144
rect -784 14123 -305 14144
rect -852 14111 -305 14123
rect -271 14111 -231 14144
rect -197 14111 -157 14144
rect -123 14136 211 14144
rect 245 14136 293 14144
rect 327 14136 375 14144
rect 409 14136 457 14144
rect 491 14136 539 14144
rect 573 14136 621 14144
rect 655 14136 703 14144
rect 737 14136 898 14144
rect -123 14111 898 14136
rect -852 14106 898 14111
rect -852 14072 -828 14106
rect -794 14085 -759 14106
rect -784 14072 -759 14085
rect -725 14072 -690 14106
rect -656 14072 -621 14106
rect -587 14072 -552 14106
rect -518 14072 -483 14106
rect -449 14072 -414 14106
rect -380 14072 -345 14106
rect -311 14073 -276 14106
rect -242 14073 -207 14106
rect -173 14073 -138 14106
rect -311 14072 -305 14073
rect -242 14072 -231 14073
rect -173 14072 -157 14073
rect -104 14072 -69 14106
rect -35 14072 0 14106
rect 34 14072 69 14106
rect 103 14072 138 14106
rect 172 14072 207 14106
rect 241 14097 276 14106
rect 310 14097 345 14106
rect 379 14097 414 14106
rect 245 14072 276 14097
rect 327 14072 345 14097
rect 409 14072 414 14097
rect 448 14097 483 14106
rect 517 14097 552 14106
rect 448 14072 457 14097
rect 517 14072 539 14097
rect 586 14072 621 14106
rect 655 14072 690 14106
rect 724 14097 759 14106
rect 737 14072 759 14097
rect 793 14072 828 14106
rect 862 14072 898 14106
rect -852 14051 -818 14072
rect -784 14051 -305 14072
rect -852 14039 -305 14051
rect -271 14039 -231 14072
rect -197 14039 -157 14072
rect -123 14063 211 14072
rect 245 14063 293 14072
rect 327 14063 375 14072
rect 409 14063 457 14072
rect 491 14063 539 14072
rect 573 14063 621 14072
rect 655 14063 703 14072
rect 737 14063 898 14072
rect -123 14039 898 14063
rect -852 14034 898 14039
rect -852 14000 -828 14034
rect -794 14013 -759 14034
rect -784 14000 -759 14013
rect -725 14000 -690 14034
rect -656 14000 -621 14034
rect -587 14000 -552 14034
rect -518 14000 -483 14034
rect -449 14000 -414 14034
rect -380 14000 -345 14034
rect -311 14001 -276 14034
rect -242 14001 -207 14034
rect -173 14001 -138 14034
rect -311 14000 -305 14001
rect -242 14000 -231 14001
rect -173 14000 -157 14001
rect -104 14000 -69 14034
rect -35 14000 0 14034
rect 34 14000 69 14034
rect 103 14000 138 14034
rect 172 14000 207 14034
rect 241 14024 276 14034
rect 310 14024 345 14034
rect 379 14024 414 14034
rect 245 14000 276 14024
rect 327 14000 345 14024
rect 409 14000 414 14024
rect 448 14024 483 14034
rect 517 14024 552 14034
rect 448 14000 457 14024
rect 517 14000 539 14024
rect 586 14000 621 14034
rect 655 14000 690 14034
rect 724 14024 759 14034
rect 737 14000 759 14024
rect 793 14000 828 14034
rect 862 14000 898 14034
rect -852 13979 -818 14000
rect -784 13979 -305 14000
rect -852 13967 -305 13979
rect -271 13967 -231 14000
rect -197 13967 -157 14000
rect -123 13996 211 14000
rect -123 13967 20 13996
rect -852 13966 20 13967
rect -852 13907 -818 13966
rect -784 13932 -748 13966
rect -714 13932 -678 13966
rect -644 13932 -608 13966
rect -574 13932 -538 13966
rect -504 13932 -468 13966
rect -434 13932 -398 13966
rect -364 13932 -328 13966
rect -294 13932 -258 13966
rect -224 13932 -188 13966
rect -154 13932 -118 13966
rect -84 13932 -48 13966
rect -14 13932 20 13966
rect -784 13929 20 13932
rect -784 13907 -305 13929
rect -852 13898 -305 13907
rect -271 13898 -231 13929
rect -197 13898 -157 13929
rect -123 13898 20 13929
rect -852 13835 -818 13898
rect -784 13864 -748 13898
rect -714 13864 -678 13898
rect -644 13864 -608 13898
rect -574 13864 -538 13898
rect -504 13864 -468 13898
rect -434 13864 -398 13898
rect -364 13864 -328 13898
rect -271 13895 -258 13898
rect -197 13895 -188 13898
rect -123 13895 -118 13898
rect -294 13864 -258 13895
rect -224 13864 -188 13895
rect -154 13864 -118 13895
rect -84 13864 -48 13898
rect -14 13864 20 13898
rect -784 13857 20 13864
rect -784 13835 -305 13857
rect -852 13830 -305 13835
rect -271 13830 -231 13857
rect -197 13830 -157 13857
rect -123 13830 20 13857
rect -852 13763 -818 13830
rect -784 13796 -748 13830
rect -714 13796 -678 13830
rect -644 13796 -608 13830
rect -574 13796 -538 13830
rect -504 13796 -468 13830
rect -434 13796 -398 13830
rect -364 13796 -328 13830
rect -271 13823 -258 13830
rect -197 13823 -188 13830
rect -123 13823 -118 13830
rect -294 13796 -258 13823
rect -224 13796 -188 13823
rect -154 13796 -118 13823
rect -84 13796 -48 13830
rect -14 13796 20 13830
rect -784 13785 20 13796
rect -784 13763 -305 13785
rect -852 13762 -305 13763
rect -271 13762 -231 13785
rect -197 13762 -157 13785
rect -123 13762 20 13785
rect -852 13728 -818 13762
rect -784 13728 -748 13762
rect -714 13728 -678 13762
rect -644 13728 -608 13762
rect -574 13728 -538 13762
rect -504 13728 -468 13762
rect -434 13728 -398 13762
rect -364 13728 -328 13762
rect -271 13751 -258 13762
rect -197 13751 -188 13762
rect -123 13751 -118 13762
rect -294 13728 -258 13751
rect -224 13728 -188 13751
rect -154 13728 -118 13751
rect -84 13728 -48 13762
rect -14 13728 20 13762
rect -852 13725 20 13728
rect -852 13660 -818 13725
rect -784 13713 20 13725
rect -784 13694 -305 13713
rect -271 13694 -231 13713
rect -197 13694 -157 13713
rect -123 13694 20 13713
rect -784 13660 -748 13694
rect -714 13660 -678 13694
rect -644 13660 -608 13694
rect -574 13660 -538 13694
rect -504 13660 -468 13694
rect -434 13660 -398 13694
rect -364 13660 -328 13694
rect -271 13679 -258 13694
rect -197 13679 -188 13694
rect -123 13679 -118 13694
rect -294 13660 -258 13679
rect -224 13660 -188 13679
rect -154 13660 -118 13679
rect -84 13660 -48 13694
rect -14 13660 20 13694
rect -852 13653 20 13660
rect -852 13592 -818 13653
rect -784 13641 20 13653
rect -784 13626 -305 13641
rect -271 13626 -231 13641
rect -197 13626 -157 13641
rect -123 13626 20 13641
rect -784 13592 -748 13626
rect -714 13592 -678 13626
rect -644 13592 -608 13626
rect -574 13592 -538 13626
rect -504 13592 -468 13626
rect -434 13592 -398 13626
rect -364 13592 -328 13626
rect -271 13607 -258 13626
rect -197 13607 -188 13626
rect -123 13607 -118 13626
rect -294 13592 -258 13607
rect -224 13592 -188 13607
rect -154 13592 -118 13607
rect -84 13592 -48 13626
rect -14 13592 20 13626
rect -852 13581 20 13592
rect -852 13524 -818 13581
rect -784 13569 20 13581
rect -784 13558 -305 13569
rect -271 13558 -231 13569
rect -197 13558 -157 13569
rect -123 13558 20 13569
rect -784 13524 -748 13558
rect -714 13524 -678 13558
rect -644 13524 -608 13558
rect -574 13524 -538 13558
rect -504 13524 -468 13558
rect -434 13524 -398 13558
rect -364 13524 -328 13558
rect -271 13535 -258 13558
rect -197 13535 -188 13558
rect -123 13535 -118 13558
rect -294 13524 -258 13535
rect -224 13524 -188 13535
rect -154 13524 -118 13535
rect -84 13524 -48 13558
rect -14 13524 20 13558
rect -852 13509 20 13524
rect -852 13456 -818 13509
rect -784 13497 20 13509
rect -784 13490 -305 13497
rect -271 13490 -231 13497
rect -197 13490 -157 13497
rect -123 13490 20 13497
rect -784 13456 -748 13490
rect -714 13456 -678 13490
rect -644 13456 -608 13490
rect -574 13456 -538 13490
rect -504 13456 -468 13490
rect -434 13456 -398 13490
rect -364 13456 -328 13490
rect -271 13463 -258 13490
rect -197 13463 -188 13490
rect -123 13463 -118 13490
rect -294 13456 -258 13463
rect -224 13456 -188 13463
rect -154 13456 -118 13463
rect -84 13456 -48 13490
rect -14 13456 20 13490
rect -852 13437 20 13456
rect -852 13388 -818 13437
rect -784 13425 20 13437
rect -784 13422 -305 13425
rect -271 13422 -231 13425
rect -197 13422 -157 13425
rect -123 13422 20 13425
rect -784 13388 -748 13422
rect -714 13388 -678 13422
rect -644 13388 -608 13422
rect -574 13388 -538 13422
rect -504 13388 -468 13422
rect -434 13388 -398 13422
rect -364 13388 -328 13422
rect -271 13391 -258 13422
rect -197 13391 -188 13422
rect -123 13391 -118 13422
rect -294 13388 -258 13391
rect -224 13388 -188 13391
rect -154 13388 -118 13391
rect -84 13388 -48 13422
rect -14 13388 20 13422
rect -852 13365 20 13388
rect -852 13320 -818 13365
rect -784 13354 20 13365
rect -784 13320 -748 13354
rect -714 13320 -678 13354
rect -644 13320 -608 13354
rect -574 13320 -538 13354
rect -504 13320 -468 13354
rect -434 13320 -398 13354
rect -364 13320 -328 13354
rect -294 13353 -258 13354
rect -224 13353 -188 13354
rect -154 13353 -118 13354
rect -271 13320 -258 13353
rect -197 13320 -188 13353
rect -123 13320 -118 13353
rect -84 13320 -48 13354
rect -14 13320 20 13354
rect -852 13319 -305 13320
rect -271 13319 -231 13320
rect -197 13319 -157 13320
rect -123 13319 20 13320
rect -852 13293 20 13319
rect -852 13252 -818 13293
rect -784 13286 20 13293
rect -784 13252 -748 13286
rect -714 13252 -678 13286
rect -644 13252 -608 13286
rect -574 13252 -538 13286
rect -504 13252 -468 13286
rect -434 13252 -398 13286
rect -364 13252 -328 13286
rect -294 13281 -258 13286
rect -224 13281 -188 13286
rect -154 13281 -118 13286
rect -271 13252 -258 13281
rect -197 13252 -188 13281
rect -123 13252 -118 13281
rect -84 13252 -48 13286
rect -14 13252 20 13286
rect -852 13247 -305 13252
rect -271 13247 -231 13252
rect -197 13247 -157 13252
rect -123 13247 20 13252
rect -852 13221 20 13247
rect -852 13184 -818 13221
rect -784 13218 20 13221
rect -784 13184 -748 13218
rect -714 13184 -678 13218
rect -644 13184 -608 13218
rect -574 13184 -538 13218
rect -504 13184 -468 13218
rect -434 13184 -398 13218
rect -364 13184 -328 13218
rect -294 13209 -258 13218
rect -224 13209 -188 13218
rect -154 13209 -118 13218
rect -271 13184 -258 13209
rect -197 13184 -188 13209
rect -123 13184 -118 13209
rect -84 13184 -48 13218
rect -14 13184 20 13218
rect -852 13175 -305 13184
rect -271 13175 -231 13184
rect -197 13175 -157 13184
rect -123 13175 20 13184
rect -852 13150 20 13175
rect -852 13115 -818 13150
rect -784 13116 -748 13150
rect -714 13116 -678 13150
rect -644 13116 -608 13150
rect -574 13116 -538 13150
rect -504 13116 -468 13150
rect -434 13116 -398 13150
rect -364 13116 -328 13150
rect -294 13137 -258 13150
rect -224 13137 -188 13150
rect -154 13137 -118 13150
rect -271 13116 -258 13137
rect -197 13116 -188 13137
rect -123 13116 -118 13137
rect -84 13116 -48 13150
rect -14 13116 20 13150
rect -784 13115 -305 13116
rect -852 13103 -305 13115
rect -271 13103 -231 13116
rect -197 13103 -157 13116
rect -123 13103 20 13116
rect -852 13082 20 13103
rect -852 13043 -818 13082
rect -784 13048 -748 13082
rect -714 13048 -678 13082
rect -644 13048 -608 13082
rect -574 13048 -538 13082
rect -504 13048 -468 13082
rect -434 13048 -398 13082
rect -364 13048 -328 13082
rect -294 13065 -258 13082
rect -224 13065 -188 13082
rect -154 13065 -118 13082
rect -271 13048 -258 13065
rect -197 13048 -188 13065
rect -123 13048 -118 13065
rect -84 13048 -48 13082
rect -14 13048 20 13082
rect -784 13043 -305 13048
rect -852 13031 -305 13043
rect -271 13031 -231 13048
rect -197 13031 -157 13048
rect -123 13031 20 13048
rect -852 13014 20 13031
rect -852 12971 -818 13014
rect -784 12980 -748 13014
rect -714 12980 -678 13014
rect -644 12980 -608 13014
rect -574 12980 -538 13014
rect -504 12980 -468 13014
rect -434 12980 -398 13014
rect -364 12980 -328 13014
rect -294 12993 -258 13014
rect -224 12993 -188 13014
rect -154 12993 -118 13014
rect -271 12980 -258 12993
rect -197 12980 -188 12993
rect -123 12980 -118 12993
rect -84 12980 -48 13014
rect -14 12980 20 13014
rect -784 12971 -305 12980
rect -852 12959 -305 12971
rect -271 12959 -231 12980
rect -197 12959 -157 12980
rect -123 12959 20 12980
rect -852 12946 20 12959
rect -852 12899 -818 12946
rect -784 12912 -748 12946
rect -714 12912 -678 12946
rect -644 12912 -608 12946
rect -574 12912 -538 12946
rect -504 12912 -468 12946
rect -434 12912 -398 12946
rect -364 12912 -328 12946
rect -294 12921 -258 12946
rect -224 12921 -188 12946
rect -154 12921 -118 12946
rect -271 12912 -258 12921
rect -197 12912 -188 12921
rect -123 12912 -118 12921
rect -84 12912 -48 12946
rect -14 12912 20 12946
rect -784 12899 -305 12912
rect -852 12887 -305 12899
rect -271 12887 -231 12912
rect -197 12887 -157 12912
rect -123 12887 20 12912
rect -852 12878 20 12887
rect -852 12827 -818 12878
rect -784 12844 -748 12878
rect -714 12844 -678 12878
rect -644 12844 -608 12878
rect -574 12844 -538 12878
rect -504 12844 -468 12878
rect -434 12844 -398 12878
rect -364 12844 -328 12878
rect -294 12849 -258 12878
rect -224 12849 -188 12878
rect -154 12849 -118 12878
rect -271 12844 -258 12849
rect -197 12844 -188 12849
rect -123 12844 -118 12849
rect -84 12844 -48 12878
rect -14 12844 20 12878
rect -784 12827 -305 12844
rect -852 12815 -305 12827
rect -271 12815 -231 12844
rect -197 12815 -157 12844
rect -123 12815 20 12844
rect -852 12810 20 12815
rect -852 12755 -818 12810
rect -784 12776 -748 12810
rect -714 12776 -678 12810
rect -644 12776 -608 12810
rect -574 12776 -538 12810
rect -504 12776 -468 12810
rect -434 12776 -398 12810
rect -364 12776 -328 12810
rect -294 12777 -258 12810
rect -224 12777 -188 12810
rect -154 12777 -118 12810
rect -271 12776 -258 12777
rect -197 12776 -188 12777
rect -123 12776 -118 12777
rect -84 12776 -48 12810
rect -14 12776 20 12810
rect -784 12755 -305 12776
rect -852 12743 -305 12755
rect -271 12743 -231 12776
rect -197 12743 -157 12776
rect -123 12743 20 12776
rect -852 12742 20 12743
rect -852 12683 -818 12742
rect -784 12708 -748 12742
rect -714 12708 -678 12742
rect -644 12708 -608 12742
rect -574 12708 -538 12742
rect -504 12708 -468 12742
rect -434 12708 -398 12742
rect -364 12708 -328 12742
rect -294 12708 -258 12742
rect -224 12708 -188 12742
rect -154 12708 -118 12742
rect -84 12708 -48 12742
rect -14 12708 20 12742
rect -784 12705 20 12708
rect -784 12683 -305 12705
rect -852 12674 -305 12683
rect -271 12674 -231 12705
rect -197 12674 -157 12705
rect -123 12674 20 12705
rect -852 12611 -818 12674
rect -784 12640 -748 12674
rect -714 12640 -678 12674
rect -644 12640 -608 12674
rect -574 12640 -538 12674
rect -504 12640 -468 12674
rect -434 12640 -398 12674
rect -364 12640 -328 12674
rect -271 12671 -258 12674
rect -197 12671 -188 12674
rect -123 12671 -118 12674
rect -294 12640 -258 12671
rect -224 12640 -188 12671
rect -154 12640 -118 12671
rect -84 12640 -48 12674
rect -14 12640 20 12674
rect -784 12633 20 12640
rect -784 12611 -305 12633
rect -852 12606 -305 12611
rect -271 12606 -231 12633
rect -197 12606 -157 12633
rect -123 12606 20 12633
rect -852 12539 -818 12606
rect -784 12572 -748 12606
rect -714 12572 -678 12606
rect -644 12572 -608 12606
rect -574 12572 -538 12606
rect -504 12572 -468 12606
rect -434 12572 -398 12606
rect -364 12572 -328 12606
rect -271 12599 -258 12606
rect -197 12599 -188 12606
rect -123 12599 -118 12606
rect -294 12572 -258 12599
rect -224 12572 -188 12599
rect -154 12572 -118 12599
rect -84 12572 -48 12606
rect -14 12572 20 12606
rect -784 12561 20 12572
rect -784 12539 -305 12561
rect -852 12538 -305 12539
rect -271 12538 -231 12561
rect -197 12538 -157 12561
rect -123 12538 20 12561
rect -852 12504 -818 12538
rect -784 12504 -748 12538
rect -714 12504 -678 12538
rect -644 12504 -608 12538
rect -574 12504 -538 12538
rect -504 12504 -468 12538
rect -434 12504 -398 12538
rect -364 12504 -328 12538
rect -271 12527 -258 12538
rect -197 12527 -188 12538
rect -123 12527 -118 12538
rect -294 12504 -258 12527
rect -224 12504 -188 12527
rect -154 12504 -118 12527
rect -84 12504 -48 12538
rect -14 12504 20 12538
rect -852 12501 20 12504
rect -852 12436 -818 12501
rect -784 12489 20 12501
rect -784 12470 -305 12489
rect -271 12470 -231 12489
rect -197 12470 -157 12489
rect -123 12470 20 12489
rect -784 12436 -748 12470
rect -714 12436 -678 12470
rect -644 12436 -608 12470
rect -574 12436 -538 12470
rect -504 12436 -468 12470
rect -434 12436 -398 12470
rect -364 12436 -328 12470
rect -271 12455 -258 12470
rect -197 12455 -188 12470
rect -123 12455 -118 12470
rect -294 12436 -258 12455
rect -224 12436 -188 12455
rect -154 12436 -118 12455
rect -84 12436 -48 12470
rect -14 12436 20 12470
rect 245 13990 293 14000
rect 327 13990 375 14000
rect 409 13990 457 14000
rect 491 13990 539 14000
rect 573 13990 621 14000
rect 655 13990 703 14000
rect 737 13996 898 14000
rect 211 13951 737 13990
rect 245 13917 293 13951
rect 327 13917 375 13951
rect 409 13917 457 13951
rect 491 13917 539 13951
rect 573 13917 621 13951
rect 655 13917 703 13951
rect 211 13878 737 13917
rect 245 13844 293 13878
rect 327 13844 375 13878
rect 409 13844 457 13878
rect 491 13844 539 13878
rect 573 13844 621 13878
rect 655 13844 703 13878
rect 211 13805 737 13844
rect 245 13771 293 13805
rect 327 13771 375 13805
rect 409 13771 457 13805
rect 491 13771 539 13805
rect 573 13771 621 13805
rect 655 13771 703 13805
rect 211 13732 737 13771
rect 245 13698 293 13732
rect 327 13698 375 13732
rect 409 13698 457 13732
rect 491 13698 539 13732
rect 573 13698 621 13732
rect 655 13698 703 13732
rect 211 13658 737 13698
rect 245 13624 293 13658
rect 327 13624 375 13658
rect 409 13624 457 13658
rect 491 13624 539 13658
rect 573 13624 621 13658
rect 655 13624 703 13658
rect 211 13584 737 13624
rect 245 13550 293 13584
rect 327 13550 375 13584
rect 409 13550 457 13584
rect 491 13550 539 13584
rect 573 13550 621 13584
rect 655 13550 703 13584
rect 211 13510 737 13550
rect 245 13476 293 13510
rect 327 13476 375 13510
rect 409 13476 457 13510
rect 491 13476 539 13510
rect 573 13476 621 13510
rect 655 13476 703 13510
rect 211 13436 737 13476
rect 245 13402 293 13436
rect 327 13402 375 13436
rect 409 13402 457 13436
rect 491 13402 539 13436
rect 573 13402 621 13436
rect 655 13402 703 13436
rect 211 13362 737 13402
rect 245 13328 293 13362
rect 327 13328 375 13362
rect 409 13328 457 13362
rect 491 13328 539 13362
rect 573 13328 621 13362
rect 655 13328 703 13362
rect 211 13288 737 13328
rect 245 13254 293 13288
rect 327 13254 375 13288
rect 409 13254 457 13288
rect 491 13254 539 13288
rect 573 13254 621 13288
rect 655 13254 703 13288
rect 211 13214 737 13254
rect 245 13180 293 13214
rect 327 13180 375 13214
rect 409 13180 457 13214
rect 491 13180 539 13214
rect 573 13180 621 13214
rect 655 13180 703 13214
rect 211 13140 737 13180
rect 245 13106 293 13140
rect 327 13106 375 13140
rect 409 13106 457 13140
rect 491 13106 539 13140
rect 573 13106 621 13140
rect 655 13106 703 13140
rect 211 13066 737 13106
rect 245 13032 293 13066
rect 327 13032 375 13066
rect 409 13032 457 13066
rect 491 13032 539 13066
rect 573 13032 621 13066
rect 655 13032 703 13066
rect 211 12992 737 13032
rect 245 12958 293 12992
rect 327 12958 375 12992
rect 409 12958 457 12992
rect 491 12958 539 12992
rect 573 12958 621 12992
rect 655 12958 703 12992
rect 211 12918 737 12958
rect 245 12884 293 12918
rect 327 12884 375 12918
rect 409 12884 457 12918
rect 491 12884 539 12918
rect 573 12884 621 12918
rect 655 12884 703 12918
rect 211 12844 737 12884
rect 245 12810 293 12844
rect 327 12810 375 12844
rect 409 12810 457 12844
rect 491 12810 539 12844
rect 573 12810 621 12844
rect 655 12810 703 12844
rect 211 12770 737 12810
rect 245 12736 293 12770
rect 327 12736 375 12770
rect 409 12736 457 12770
rect 491 12736 539 12770
rect 573 12736 621 12770
rect 655 12736 703 12770
rect 211 12696 737 12736
rect 245 12662 293 12696
rect 327 12662 375 12696
rect 409 12662 457 12696
rect 491 12662 539 12696
rect 573 12662 621 12696
rect 655 12662 703 12696
rect 211 12622 737 12662
rect 245 12588 293 12622
rect 327 12588 375 12622
rect 409 12588 457 12622
rect 491 12588 539 12622
rect 573 12588 621 12622
rect 655 12588 703 12622
rect 211 12548 737 12588
rect 245 12514 293 12548
rect 327 12514 375 12548
rect 409 12514 457 12548
rect 491 12514 539 12548
rect 573 12514 621 12548
rect 655 12514 703 12548
rect 211 12474 737 12514
rect 245 12440 293 12474
rect 327 12440 375 12474
rect 409 12440 457 12474
rect 491 12440 539 12474
rect 573 12440 621 12474
rect 655 12440 703 12474
rect -852 12429 20 12436
rect -852 12368 -818 12429
rect -784 12417 20 12429
rect -784 12402 -305 12417
rect -271 12402 -231 12417
rect -197 12402 -157 12417
rect -123 12402 20 12417
rect -784 12368 -748 12402
rect -714 12368 -678 12402
rect -644 12368 -608 12402
rect -574 12368 -538 12402
rect -504 12368 -468 12402
rect -434 12368 -398 12402
rect -364 12368 -328 12402
rect -271 12383 -258 12402
rect -197 12383 -188 12402
rect -123 12383 -118 12402
rect -294 12368 -258 12383
rect -224 12368 -188 12383
rect -154 12368 -118 12383
rect -84 12368 -48 12402
rect -14 12368 20 12402
rect -852 12357 20 12368
rect -852 12300 -818 12357
rect -784 12345 20 12357
rect -784 12334 -305 12345
rect -271 12334 -231 12345
rect -197 12334 -157 12345
rect -123 12334 20 12345
rect -784 12300 -748 12334
rect -714 12300 -678 12334
rect -644 12300 -608 12334
rect -574 12300 -538 12334
rect -504 12300 -468 12334
rect -434 12300 -398 12334
rect -364 12300 -328 12334
rect -271 12311 -258 12334
rect -197 12311 -188 12334
rect -123 12311 -118 12334
rect -294 12300 -258 12311
rect -224 12300 -188 12311
rect -154 12300 -118 12311
rect -84 12300 -48 12334
rect -14 12300 20 12334
rect -852 12285 20 12300
rect -852 12232 -818 12285
rect -784 12273 20 12285
rect -784 12266 -305 12273
rect -271 12266 -231 12273
rect -197 12266 -157 12273
rect -123 12266 20 12273
rect -784 12232 -748 12266
rect -714 12232 -678 12266
rect -644 12232 -608 12266
rect -574 12232 -538 12266
rect -504 12232 -468 12266
rect -434 12232 -398 12266
rect -364 12232 -328 12266
rect -271 12239 -258 12266
rect -197 12239 -188 12266
rect -123 12239 -118 12266
rect -294 12232 -258 12239
rect -224 12232 -188 12239
rect -154 12232 -118 12239
rect -84 12232 -48 12266
rect -14 12232 20 12266
rect -852 12213 20 12232
rect -852 12164 -818 12213
rect -784 12201 20 12213
rect -784 12198 -305 12201
rect -271 12198 -231 12201
rect -197 12198 -157 12201
rect -123 12198 20 12201
rect -784 12164 -748 12198
rect -714 12164 -678 12198
rect -644 12164 -608 12198
rect -574 12164 -538 12198
rect -504 12164 -468 12198
rect -434 12164 -398 12198
rect -364 12164 -328 12198
rect -271 12167 -258 12198
rect -197 12167 -188 12198
rect -123 12167 -118 12198
rect -294 12164 -258 12167
rect -224 12164 -188 12167
rect -154 12164 -118 12167
rect -84 12164 -48 12198
rect -14 12164 20 12198
rect -852 12160 20 12164
rect -852 12141 68 12160
rect -852 12096 -818 12141
rect -784 12130 68 12141
rect -784 12096 -748 12130
rect -714 12096 -678 12130
rect -644 12096 -608 12130
rect -574 12096 -538 12130
rect -504 12096 -468 12130
rect -434 12096 -398 12130
rect -364 12096 -328 12130
rect -294 12129 -258 12130
rect -224 12129 -188 12130
rect -154 12129 -118 12130
rect -271 12096 -258 12129
rect -197 12096 -188 12129
rect -123 12096 -118 12129
rect -84 12096 -48 12130
rect -14 12096 68 12130
rect -852 12095 -305 12096
rect -271 12095 -231 12096
rect -197 12095 -157 12096
rect -123 12095 68 12096
rect -852 12069 68 12095
rect -852 12028 -818 12069
rect -784 12062 68 12069
rect -784 12028 -748 12062
rect -714 12028 -678 12062
rect -644 12028 -608 12062
rect -574 12028 -538 12062
rect -504 12028 -468 12062
rect -434 12028 -398 12062
rect -364 12028 -328 12062
rect -294 12057 -258 12062
rect -224 12057 -188 12062
rect -154 12057 -118 12062
rect -271 12028 -258 12057
rect -197 12028 -188 12057
rect -123 12028 -118 12057
rect -84 12028 -48 12062
rect -14 12028 68 12062
rect -852 12023 -305 12028
rect -271 12023 -231 12028
rect -197 12023 -157 12028
rect -123 12023 68 12028
rect -852 11997 68 12023
rect -852 11960 -818 11997
rect -784 11994 68 11997
rect -784 11960 -748 11994
rect -714 11960 -678 11994
rect -644 11960 -608 11994
rect -574 11960 -538 11994
rect -504 11960 -468 11994
rect -434 11960 -398 11994
rect -364 11960 -328 11994
rect -294 11985 -258 11994
rect -224 11985 -188 11994
rect -154 11985 -118 11994
rect -271 11960 -258 11985
rect -197 11960 -188 11985
rect -123 11960 -118 11985
rect -84 11960 -48 11994
rect -14 11960 68 11994
rect -852 11951 -305 11960
rect -271 11951 -231 11960
rect -197 11951 -157 11960
rect -123 11951 68 11960
rect -852 11926 68 11951
rect -852 11891 -818 11926
rect -784 11892 -748 11926
rect -714 11892 -678 11926
rect -644 11892 -608 11926
rect -574 11892 -538 11926
rect -504 11892 -468 11926
rect -434 11892 -398 11926
rect -364 11892 -328 11926
rect -294 11913 -258 11926
rect -224 11913 -188 11926
rect -154 11913 -118 11926
rect -271 11892 -258 11913
rect -197 11892 -188 11913
rect -123 11892 -118 11913
rect -84 11892 -48 11926
rect -14 11892 68 11926
rect -784 11891 -305 11892
rect -852 11879 -305 11891
rect -271 11879 -231 11892
rect -197 11879 -157 11892
rect -123 11879 68 11892
rect -852 11858 68 11879
rect -852 11819 -818 11858
rect -784 11824 -748 11858
rect -714 11824 -678 11858
rect -644 11824 -608 11858
rect -574 11824 -538 11858
rect -504 11824 -468 11858
rect -434 11824 -398 11858
rect -364 11824 -328 11858
rect -294 11841 -258 11858
rect -224 11841 -188 11858
rect -154 11841 -118 11858
rect -271 11824 -258 11841
rect -197 11824 -188 11841
rect -123 11824 -118 11841
rect -84 11824 -48 11858
rect -14 11824 68 11858
rect -784 11819 -305 11824
rect -852 11807 -305 11819
rect -271 11807 -231 11824
rect -197 11807 -157 11824
rect -123 11807 68 11824
rect -852 11790 68 11807
rect -852 11747 -818 11790
rect -784 11756 -748 11790
rect -714 11756 -678 11790
rect -644 11756 -608 11790
rect -574 11756 -538 11790
rect -504 11756 -468 11790
rect -434 11756 -398 11790
rect -364 11756 -328 11790
rect -294 11769 -258 11790
rect -224 11769 -188 11790
rect -154 11769 -118 11790
rect -271 11756 -258 11769
rect -197 11756 -188 11769
rect -123 11756 -118 11769
rect -84 11756 -48 11790
rect -14 11756 68 11790
rect -784 11747 -305 11756
rect -852 11735 -305 11747
rect -271 11735 -231 11756
rect -197 11735 -157 11756
rect -123 11735 68 11756
rect -852 11722 68 11735
rect -852 11675 -818 11722
rect -784 11688 -748 11722
rect -714 11688 -678 11722
rect -644 11688 -608 11722
rect -574 11688 -538 11722
rect -504 11688 -468 11722
rect -434 11688 -398 11722
rect -364 11688 -328 11722
rect -294 11697 -258 11722
rect -224 11697 -188 11722
rect -154 11697 -118 11722
rect -271 11688 -258 11697
rect -197 11688 -188 11697
rect -123 11688 -118 11697
rect -84 11688 -48 11722
rect -14 11688 68 11722
rect -784 11675 -305 11688
rect -852 11663 -305 11675
rect -271 11663 -231 11688
rect -197 11663 -157 11688
rect -123 11663 68 11688
rect -852 11654 68 11663
rect -852 11603 -818 11654
rect -784 11620 -748 11654
rect -714 11620 -678 11654
rect -644 11620 -608 11654
rect -574 11620 -538 11654
rect -504 11620 -468 11654
rect -434 11620 -398 11654
rect -364 11620 -328 11654
rect -294 11625 -258 11654
rect -224 11625 -188 11654
rect -154 11625 -118 11654
rect -271 11620 -258 11625
rect -197 11620 -188 11625
rect -123 11620 -118 11625
rect -84 11620 -48 11654
rect -14 11620 68 11654
rect -784 11603 -305 11620
rect -852 11591 -305 11603
rect -271 11591 -231 11620
rect -197 11591 -157 11620
rect -123 11591 68 11620
rect -852 11586 68 11591
rect -852 11531 -818 11586
rect -784 11552 -748 11586
rect -714 11552 -678 11586
rect -644 11552 -608 11586
rect -574 11552 -538 11586
rect -504 11552 -468 11586
rect -434 11552 -398 11586
rect -364 11552 -328 11586
rect -294 11553 -258 11586
rect -224 11553 -188 11586
rect -154 11553 -118 11586
rect -271 11552 -258 11553
rect -197 11552 -188 11553
rect -123 11552 -118 11553
rect -84 11552 -48 11586
rect -14 11552 68 11586
rect -784 11531 -305 11552
rect -852 11519 -305 11531
rect -271 11519 -231 11552
rect -197 11519 -157 11552
rect -123 11519 68 11552
rect -852 11518 68 11519
rect -852 11459 -818 11518
rect -784 11484 -748 11518
rect -714 11484 -678 11518
rect -644 11484 -608 11518
rect -574 11484 -538 11518
rect -504 11484 -468 11518
rect -434 11484 -398 11518
rect -364 11484 -328 11518
rect -294 11484 -258 11518
rect -224 11484 -188 11518
rect -154 11484 -118 11518
rect -84 11484 -48 11518
rect -14 11484 68 11518
rect -784 11481 68 11484
rect -784 11459 -305 11481
rect -852 11450 -305 11459
rect -271 11450 -231 11481
rect -197 11450 -157 11481
rect -123 11450 68 11481
rect -852 11387 -818 11450
rect -784 11416 -748 11450
rect -714 11416 -678 11450
rect -644 11416 -608 11450
rect -574 11416 -538 11450
rect -504 11416 -468 11450
rect -434 11416 -398 11450
rect -364 11416 -328 11450
rect -271 11447 -258 11450
rect -197 11447 -188 11450
rect -123 11447 -118 11450
rect -294 11416 -258 11447
rect -224 11416 -188 11447
rect -154 11416 -118 11447
rect -84 11416 -48 11450
rect -14 11416 68 11450
rect -784 11409 68 11416
rect -784 11387 -305 11409
rect -852 11382 -305 11387
rect -271 11382 -231 11409
rect -197 11382 -157 11409
rect -123 11382 68 11409
rect -852 11315 -818 11382
rect -784 11348 -748 11382
rect -714 11348 -678 11382
rect -644 11348 -608 11382
rect -574 11348 -538 11382
rect -504 11348 -468 11382
rect -434 11348 -398 11382
rect -364 11348 -328 11382
rect -271 11375 -258 11382
rect -197 11375 -188 11382
rect -123 11375 -118 11382
rect -294 11348 -258 11375
rect -224 11348 -188 11375
rect -154 11348 -118 11375
rect -84 11348 -48 11382
rect -14 11348 68 11382
rect -784 11337 68 11348
rect -784 11315 -305 11337
rect -852 11314 -305 11315
rect -271 11314 -231 11337
rect -197 11314 -157 11337
rect -123 11314 68 11337
rect -852 11280 -818 11314
rect -784 11280 -748 11314
rect -714 11280 -678 11314
rect -644 11280 -608 11314
rect -574 11280 -538 11314
rect -504 11280 -468 11314
rect -434 11280 -398 11314
rect -364 11280 -328 11314
rect -271 11303 -258 11314
rect -197 11303 -188 11314
rect -123 11303 -118 11314
rect -294 11280 -258 11303
rect -224 11280 -188 11303
rect -154 11280 -118 11303
rect -84 11280 -48 11314
rect -14 11280 68 11314
rect -852 11277 68 11280
rect -852 11212 -818 11277
rect -784 11265 68 11277
rect -784 11246 -305 11265
rect -271 11246 -231 11265
rect -197 11246 -157 11265
rect -123 11246 68 11265
rect -784 11212 -748 11246
rect -714 11212 -678 11246
rect -644 11212 -608 11246
rect -574 11212 -538 11246
rect -504 11212 -468 11246
rect -434 11212 -398 11246
rect -364 11212 -328 11246
rect -271 11231 -258 11246
rect -197 11231 -188 11246
rect -123 11231 -118 11246
rect -294 11212 -258 11231
rect -224 11212 -188 11231
rect -154 11212 -118 11231
rect -84 11212 -48 11246
rect -14 11212 68 11246
rect -852 11205 68 11212
rect -852 11144 -818 11205
rect -784 11193 68 11205
rect -784 11178 -305 11193
rect -271 11178 -231 11193
rect -197 11178 -157 11193
rect -123 11178 68 11193
rect -784 11144 -748 11178
rect -714 11144 -678 11178
rect -644 11144 -608 11178
rect -574 11144 -538 11178
rect -504 11144 -468 11178
rect -434 11144 -398 11178
rect -364 11144 -328 11178
rect -271 11159 -258 11178
rect -197 11159 -188 11178
rect -123 11159 -118 11178
rect -294 11144 -258 11159
rect -224 11144 -188 11159
rect -154 11144 -118 11159
rect -84 11144 -48 11178
rect -14 11144 68 11178
rect -852 11133 68 11144
rect -852 11076 -818 11133
rect -784 11121 68 11133
rect -784 11110 -305 11121
rect -271 11110 -231 11121
rect -197 11110 -157 11121
rect -123 11110 68 11121
rect -784 11076 -748 11110
rect -714 11076 -678 11110
rect -644 11076 -608 11110
rect -574 11076 -538 11110
rect -504 11076 -468 11110
rect -434 11076 -398 11110
rect -364 11076 -328 11110
rect -271 11087 -258 11110
rect -197 11087 -188 11110
rect -123 11087 -118 11110
rect -294 11076 -258 11087
rect -224 11076 -188 11087
rect -154 11076 -118 11087
rect -84 11076 -48 11110
rect -14 11076 68 11110
rect -852 11061 68 11076
rect -852 11008 -818 11061
rect -784 11049 68 11061
rect -784 11042 -305 11049
rect -271 11042 -231 11049
rect -197 11042 -157 11049
rect -123 11042 68 11049
rect -784 11008 -748 11042
rect -714 11008 -678 11042
rect -644 11008 -608 11042
rect -574 11008 -538 11042
rect -504 11008 -468 11042
rect -434 11008 -398 11042
rect -364 11008 -328 11042
rect -271 11015 -258 11042
rect -197 11015 -188 11042
rect -123 11015 -118 11042
rect -294 11008 -258 11015
rect -224 11008 -188 11015
rect -154 11008 -118 11015
rect -84 11008 -48 11042
rect -14 11008 68 11042
rect -852 10989 68 11008
rect -852 10940 -818 10989
rect -784 10977 68 10989
rect -784 10974 -305 10977
rect -271 10974 -231 10977
rect -197 10974 -157 10977
rect -123 10974 68 10977
rect -784 10940 -748 10974
rect -714 10940 -678 10974
rect -644 10940 -608 10974
rect -574 10940 -538 10974
rect -504 10940 -468 10974
rect -434 10940 -398 10974
rect -364 10940 -328 10974
rect -271 10943 -258 10974
rect -197 10943 -188 10974
rect -123 10943 -118 10974
rect -294 10940 -258 10943
rect -224 10940 -188 10943
rect -154 10940 -118 10943
rect -84 10940 -48 10974
rect -14 10940 68 10974
rect -852 10917 68 10940
rect -852 10872 -818 10917
rect -784 10906 68 10917
rect -784 10872 -748 10906
rect -714 10872 -678 10906
rect -644 10872 -608 10906
rect -574 10872 -538 10906
rect -504 10872 -468 10906
rect -434 10872 -398 10906
rect -364 10872 -328 10906
rect -294 10905 -258 10906
rect -224 10905 -188 10906
rect -154 10905 -118 10906
rect -271 10872 -258 10905
rect -197 10872 -188 10905
rect -123 10872 -118 10905
rect -84 10872 -48 10906
rect -14 10872 68 10906
rect -852 10871 -305 10872
rect -271 10871 -231 10872
rect -197 10871 -157 10872
rect -123 10871 68 10872
rect -852 10845 68 10871
rect -852 10804 -818 10845
rect -784 10838 68 10845
rect -784 10804 -748 10838
rect -714 10804 -678 10838
rect -644 10804 -608 10838
rect -574 10804 -538 10838
rect -504 10804 -468 10838
rect -434 10804 -398 10838
rect -364 10804 -328 10838
rect -294 10833 -258 10838
rect -224 10833 -188 10838
rect -154 10833 -118 10838
rect -271 10804 -258 10833
rect -197 10804 -188 10833
rect -123 10804 -118 10833
rect -84 10804 -48 10838
rect -14 10804 68 10838
rect -852 10799 -305 10804
rect -271 10799 -231 10804
rect -197 10799 -157 10804
rect -123 10799 68 10804
rect -852 10773 68 10799
rect -852 10736 -818 10773
rect -784 10770 68 10773
rect -784 10736 -748 10770
rect -714 10736 -678 10770
rect -644 10736 -608 10770
rect -574 10736 -538 10770
rect -504 10736 -468 10770
rect -434 10736 -398 10770
rect -364 10736 -328 10770
rect -294 10761 -258 10770
rect -224 10761 -188 10770
rect -154 10761 -118 10770
rect -271 10736 -258 10761
rect -197 10736 -188 10761
rect -123 10736 -118 10761
rect -84 10736 -48 10770
rect -14 10736 68 10770
rect -852 10727 -305 10736
rect -271 10727 -231 10736
rect -197 10727 -157 10736
rect -123 10727 68 10736
rect -852 10702 68 10727
rect -852 10667 -818 10702
rect -784 10668 -748 10702
rect -714 10668 -678 10702
rect -644 10668 -608 10702
rect -574 10668 -538 10702
rect -504 10668 -468 10702
rect -434 10668 -398 10702
rect -364 10668 -328 10702
rect -294 10689 -258 10702
rect -224 10689 -188 10702
rect -154 10689 -118 10702
rect -271 10668 -258 10689
rect -197 10668 -188 10689
rect -123 10668 -118 10689
rect -84 10668 -48 10702
rect -14 10668 68 10702
rect -784 10667 -305 10668
rect -852 10655 -305 10667
rect -271 10655 -231 10668
rect -197 10655 -157 10668
rect -123 10655 68 10668
rect -852 10634 68 10655
rect -852 10595 -818 10634
rect -784 10600 -748 10634
rect -714 10600 -678 10634
rect -644 10600 -608 10634
rect -574 10600 -538 10634
rect -504 10600 -468 10634
rect -434 10600 -398 10634
rect -364 10600 -328 10634
rect -294 10617 -258 10634
rect -224 10617 -188 10634
rect -154 10617 -118 10634
rect -271 10600 -258 10617
rect -197 10600 -188 10617
rect -123 10600 -118 10617
rect -84 10600 -48 10634
rect -14 10600 68 10634
rect -784 10595 -305 10600
rect -852 10583 -305 10595
rect -271 10583 -231 10600
rect -197 10583 -157 10600
rect -123 10583 68 10600
rect -852 10566 68 10583
rect -852 10523 -818 10566
rect -784 10532 -748 10566
rect -714 10532 -678 10566
rect -644 10532 -608 10566
rect -574 10532 -538 10566
rect -504 10532 -468 10566
rect -434 10532 -398 10566
rect -364 10532 -328 10566
rect -294 10545 -258 10566
rect -224 10545 -188 10566
rect -154 10545 -118 10566
rect -271 10532 -258 10545
rect -197 10532 -188 10545
rect -123 10532 -118 10545
rect -84 10532 -48 10566
rect -14 10532 68 10566
rect -784 10523 -305 10532
rect -852 10511 -305 10523
rect -271 10511 -231 10532
rect -197 10511 -157 10532
rect -123 10511 68 10532
rect -852 10498 68 10511
rect -852 10451 -818 10498
rect -784 10464 -748 10498
rect -714 10464 -678 10498
rect -644 10464 -608 10498
rect -574 10464 -538 10498
rect -504 10464 -468 10498
rect -434 10464 -398 10498
rect -364 10464 -328 10498
rect -294 10473 -258 10498
rect -224 10473 -188 10498
rect -154 10473 -118 10498
rect -271 10464 -258 10473
rect -197 10464 -188 10473
rect -123 10464 -118 10473
rect -84 10464 -48 10498
rect -14 10464 68 10498
rect -784 10451 -305 10464
rect -852 10439 -305 10451
rect -271 10439 -231 10464
rect -197 10439 -157 10464
rect -123 10439 68 10464
rect -852 10430 68 10439
rect -852 10379 -818 10430
rect -784 10396 -748 10430
rect -714 10396 -678 10430
rect -644 10396 -608 10430
rect -574 10396 -538 10430
rect -504 10396 -468 10430
rect -434 10396 -398 10430
rect -364 10396 -328 10430
rect -294 10401 -258 10430
rect -224 10401 -188 10430
rect -154 10401 -118 10430
rect -271 10396 -258 10401
rect -197 10396 -188 10401
rect -123 10396 -118 10401
rect -84 10396 -48 10430
rect -14 10396 68 10430
rect -784 10379 -305 10396
rect -852 10367 -305 10379
rect -271 10367 -231 10396
rect -197 10367 -157 10396
rect -123 10367 68 10396
rect -852 10362 68 10367
rect -852 10307 -818 10362
rect -784 10328 -748 10362
rect -714 10328 -678 10362
rect -644 10328 -608 10362
rect -574 10328 -538 10362
rect -504 10328 -468 10362
rect -434 10328 -398 10362
rect -364 10328 -328 10362
rect -294 10329 -258 10362
rect -224 10329 -188 10362
rect -154 10329 -118 10362
rect -271 10328 -258 10329
rect -197 10328 -188 10329
rect -123 10328 -118 10329
rect -84 10328 -48 10362
rect -14 10328 68 10362
rect -784 10307 -305 10328
rect -852 10295 -305 10307
rect -271 10295 -231 10328
rect -197 10295 -157 10328
rect -123 10295 68 10328
rect -852 10294 68 10295
rect -852 10235 -818 10294
rect -784 10260 -748 10294
rect -714 10260 -678 10294
rect -644 10260 -608 10294
rect -574 10260 -538 10294
rect -504 10260 -468 10294
rect -434 10260 -398 10294
rect -364 10260 -328 10294
rect -294 10260 -258 10294
rect -224 10260 -188 10294
rect -154 10260 -118 10294
rect -84 10260 -48 10294
rect -14 10260 68 10294
rect -784 10257 68 10260
rect -784 10235 -305 10257
rect -852 10226 -305 10235
rect -271 10226 -231 10257
rect -197 10226 -157 10257
rect -123 10226 68 10257
rect -852 10163 -818 10226
rect -784 10192 -748 10226
rect -714 10192 -678 10226
rect -644 10192 -608 10226
rect -574 10192 -538 10226
rect -504 10192 -468 10226
rect -434 10192 -398 10226
rect -364 10192 -328 10226
rect -271 10223 -258 10226
rect -197 10223 -188 10226
rect -123 10223 -118 10226
rect -294 10192 -258 10223
rect -224 10192 -188 10223
rect -154 10192 -118 10223
rect -84 10192 -48 10226
rect -14 10192 68 10226
rect -784 10185 68 10192
rect -784 10163 -305 10185
rect -852 10158 -305 10163
rect -271 10158 -231 10185
rect -197 10158 -157 10185
rect -123 10158 68 10185
rect -852 10091 -818 10158
rect -784 10124 -748 10158
rect -714 10124 -678 10158
rect -644 10124 -608 10158
rect -574 10124 -538 10158
rect -504 10124 -468 10158
rect -434 10124 -398 10158
rect -364 10124 -328 10158
rect -271 10151 -258 10158
rect -197 10151 -188 10158
rect -123 10151 -118 10158
rect -294 10124 -258 10151
rect -224 10124 -188 10151
rect -154 10124 -118 10151
rect -84 10124 -48 10158
rect -14 10124 68 10158
rect -784 10113 68 10124
rect -784 10091 -305 10113
rect -852 10090 -305 10091
rect -271 10090 -231 10113
rect -197 10090 -157 10113
rect -123 10090 68 10113
rect -852 10056 -818 10090
rect -784 10056 -748 10090
rect -714 10056 -678 10090
rect -644 10056 -608 10090
rect -574 10056 -538 10090
rect -504 10056 -468 10090
rect -434 10056 -398 10090
rect -364 10056 -328 10090
rect -271 10079 -258 10090
rect -197 10079 -188 10090
rect -123 10079 -118 10090
rect -294 10056 -258 10079
rect -224 10056 -188 10079
rect -154 10056 -118 10079
rect -84 10056 -48 10090
rect -14 10056 68 10090
rect -852 10053 68 10056
rect -852 9988 -818 10053
rect -784 10041 68 10053
rect -784 10022 -305 10041
rect -271 10022 -231 10041
rect -197 10022 -157 10041
rect -123 10022 68 10041
rect -784 9988 -748 10022
rect -714 9988 -678 10022
rect -644 9988 -608 10022
rect -574 9988 -538 10022
rect -504 9988 -468 10022
rect -434 9988 -398 10022
rect -364 9988 -328 10022
rect -271 10007 -258 10022
rect -197 10007 -188 10022
rect -123 10007 -118 10022
rect -294 9988 -258 10007
rect -224 9988 -188 10007
rect -154 9988 -118 10007
rect -84 9988 -48 10022
rect -14 9988 68 10022
rect -852 9981 68 9988
rect -852 9920 -818 9981
rect -784 9969 68 9981
rect -784 9954 -305 9969
rect -271 9954 -231 9969
rect -197 9954 -157 9969
rect -123 9954 68 9969
rect -784 9920 -748 9954
rect -714 9920 -678 9954
rect -644 9920 -608 9954
rect -574 9920 -538 9954
rect -504 9920 -468 9954
rect -434 9920 -398 9954
rect -364 9920 -328 9954
rect -271 9935 -258 9954
rect -197 9935 -188 9954
rect -123 9935 -118 9954
rect -294 9920 -258 9935
rect -224 9920 -188 9935
rect -154 9920 -118 9935
rect -84 9920 -48 9954
rect -14 9920 68 9954
rect -852 9909 68 9920
rect -852 9852 -818 9909
rect -784 9897 68 9909
rect -784 9886 -305 9897
rect -271 9886 -231 9897
rect -197 9886 -157 9897
rect -123 9886 68 9897
rect -784 9852 -748 9886
rect -714 9852 -678 9886
rect -644 9852 -608 9886
rect -574 9852 -538 9886
rect -504 9852 -468 9886
rect -434 9852 -398 9886
rect -364 9852 -328 9886
rect -271 9863 -258 9886
rect -197 9863 -188 9886
rect -123 9863 -118 9886
rect -294 9852 -258 9863
rect -224 9852 -188 9863
rect -154 9852 -118 9863
rect -84 9852 -48 9886
rect -14 9852 68 9886
rect -852 9837 68 9852
rect -852 9784 -818 9837
rect -784 9825 68 9837
rect -784 9818 -305 9825
rect -271 9818 -231 9825
rect -197 9818 -157 9825
rect -123 9818 68 9825
rect -784 9784 -748 9818
rect -714 9784 -678 9818
rect -644 9784 -608 9818
rect -574 9784 -538 9818
rect -504 9784 -468 9818
rect -434 9784 -398 9818
rect -364 9784 -328 9818
rect -271 9791 -258 9818
rect -197 9791 -188 9818
rect -123 9791 -118 9818
rect -294 9784 -258 9791
rect -224 9784 -188 9791
rect -154 9784 -118 9791
rect -84 9784 -48 9818
rect -14 9784 68 9818
rect -852 9765 68 9784
rect -852 9716 -818 9765
rect -784 9753 68 9765
rect -784 9750 -305 9753
rect -271 9750 -231 9753
rect -197 9750 -157 9753
rect -123 9750 68 9753
rect -784 9716 -748 9750
rect -714 9716 -678 9750
rect -644 9716 -608 9750
rect -574 9716 -538 9750
rect -504 9716 -468 9750
rect -434 9716 -398 9750
rect -364 9716 -328 9750
rect -271 9719 -258 9750
rect -197 9719 -188 9750
rect -123 9719 -118 9750
rect -294 9716 -258 9719
rect -224 9716 -188 9719
rect -154 9716 -118 9719
rect -84 9716 -48 9750
rect -14 9716 68 9750
rect -852 9693 68 9716
rect -852 9648 -818 9693
rect -784 9682 68 9693
rect -784 9648 -748 9682
rect -714 9648 -678 9682
rect -644 9648 -608 9682
rect -574 9648 -538 9682
rect -504 9648 -468 9682
rect -434 9648 -398 9682
rect -364 9648 -328 9682
rect -294 9681 -258 9682
rect -224 9681 -188 9682
rect -154 9681 -118 9682
rect -271 9648 -258 9681
rect -197 9648 -188 9681
rect -123 9648 -118 9681
rect -84 9648 -48 9682
rect -14 9648 68 9682
rect -852 9647 -305 9648
rect -271 9647 -231 9648
rect -197 9647 -157 9648
rect -123 9647 68 9648
rect -852 9621 68 9647
rect -852 9580 -818 9621
rect -784 9614 68 9621
rect -784 9580 -748 9614
rect -714 9580 -678 9614
rect -644 9580 -608 9614
rect -574 9580 -538 9614
rect -504 9580 -468 9614
rect -434 9580 -398 9614
rect -364 9580 -328 9614
rect -294 9609 -258 9614
rect -224 9609 -188 9614
rect -154 9609 -118 9614
rect -271 9580 -258 9609
rect -197 9580 -188 9609
rect -123 9580 -118 9609
rect -84 9580 -48 9614
rect -14 9580 68 9614
rect -852 9575 -305 9580
rect -271 9575 -231 9580
rect -197 9575 -157 9580
rect -123 9575 68 9580
rect -852 9549 68 9575
rect -852 9512 -818 9549
rect -784 9546 68 9549
rect -784 9512 -748 9546
rect -714 9512 -678 9546
rect -644 9512 -608 9546
rect -574 9512 -538 9546
rect -504 9512 -468 9546
rect -434 9512 -398 9546
rect -364 9512 -328 9546
rect -294 9537 -258 9546
rect -224 9537 -188 9546
rect -154 9537 -118 9546
rect -271 9512 -258 9537
rect -197 9512 -188 9537
rect -123 9512 -118 9537
rect -84 9512 -48 9546
rect -14 9512 68 9546
rect -852 9503 -305 9512
rect -271 9503 -231 9512
rect -197 9503 -157 9512
rect -123 9503 68 9512
rect -852 9478 68 9503
rect -852 9443 -818 9478
rect -784 9444 -748 9478
rect -714 9444 -678 9478
rect -644 9444 -608 9478
rect -574 9444 -538 9478
rect -504 9444 -468 9478
rect -434 9444 -398 9478
rect -364 9444 -328 9478
rect -294 9465 -258 9478
rect -224 9465 -188 9478
rect -154 9465 -118 9478
rect -271 9444 -258 9465
rect -197 9444 -188 9465
rect -123 9444 -118 9465
rect -84 9444 -48 9478
rect -14 9444 68 9478
rect -784 9443 -305 9444
rect -852 9431 -305 9443
rect -271 9431 -231 9444
rect -197 9431 -157 9444
rect -123 9431 68 9444
rect -852 9410 68 9431
rect -852 9371 -818 9410
rect -784 9376 -748 9410
rect -714 9376 -678 9410
rect -644 9376 -608 9410
rect -574 9376 -538 9410
rect -504 9376 -468 9410
rect -434 9376 -398 9410
rect -364 9376 -328 9410
rect -294 9393 -258 9410
rect -224 9393 -188 9410
rect -154 9393 -118 9410
rect -271 9376 -258 9393
rect -197 9376 -188 9393
rect -123 9376 -118 9393
rect -84 9376 -48 9410
rect -14 9376 68 9410
rect -784 9371 -305 9376
rect -852 9359 -305 9371
rect -271 9359 -231 9376
rect -197 9359 -157 9376
rect -123 9359 68 9376
rect -852 9342 68 9359
rect -852 9299 -818 9342
rect -784 9308 -748 9342
rect -714 9308 -678 9342
rect -644 9308 -608 9342
rect -574 9308 -538 9342
rect -504 9308 -468 9342
rect -434 9308 -398 9342
rect -364 9308 -328 9342
rect -294 9321 -258 9342
rect -224 9321 -188 9342
rect -154 9321 -118 9342
rect -271 9308 -258 9321
rect -197 9308 -188 9321
rect -123 9308 -118 9321
rect -84 9308 -48 9342
rect -14 9308 68 9342
rect -784 9299 -305 9308
rect -852 9287 -305 9299
rect -271 9287 -231 9308
rect -197 9287 -157 9308
rect -123 9287 68 9308
rect -852 9274 68 9287
rect -852 9227 -818 9274
rect -784 9240 -748 9274
rect -714 9240 -678 9274
rect -644 9240 -608 9274
rect -574 9240 -538 9274
rect -504 9240 -468 9274
rect -434 9240 -398 9274
rect -364 9240 -328 9274
rect -294 9249 -258 9274
rect -224 9249 -188 9274
rect -154 9249 -118 9274
rect -271 9240 -258 9249
rect -197 9240 -188 9249
rect -123 9240 -118 9249
rect -84 9240 -48 9274
rect -14 9240 68 9274
rect -784 9227 -305 9240
rect -852 9215 -305 9227
rect -271 9215 -231 9240
rect -197 9215 -157 9240
rect -123 9215 68 9240
rect -852 9206 68 9215
rect -852 9155 -818 9206
rect -784 9172 -748 9206
rect -714 9172 -678 9206
rect -644 9172 -608 9206
rect -574 9172 -538 9206
rect -504 9172 -468 9206
rect -434 9172 -398 9206
rect -364 9172 -328 9206
rect -294 9177 -258 9206
rect -224 9177 -188 9206
rect -154 9177 -118 9206
rect -271 9172 -258 9177
rect -197 9172 -188 9177
rect -123 9172 -118 9177
rect -84 9172 -48 9206
rect -14 9172 68 9206
rect -784 9155 -305 9172
rect -852 9143 -305 9155
rect -271 9143 -231 9172
rect -197 9143 -157 9172
rect -123 9143 68 9172
rect -852 9138 68 9143
rect -852 9083 -818 9138
rect -784 9104 -748 9138
rect -714 9104 -678 9138
rect -644 9104 -608 9138
rect -574 9104 -538 9138
rect -504 9104 -468 9138
rect -434 9104 -398 9138
rect -364 9104 -328 9138
rect -294 9105 -258 9138
rect -224 9105 -188 9138
rect -154 9105 -118 9138
rect -271 9104 -258 9105
rect -197 9104 -188 9105
rect -123 9104 -118 9105
rect -84 9104 -48 9138
rect -14 9104 68 9138
rect -784 9083 -305 9104
rect -852 9071 -305 9083
rect -271 9071 -231 9104
rect -197 9071 -157 9104
rect -123 9071 68 9104
rect -852 9070 68 9071
rect -852 9011 -818 9070
rect -784 9036 -748 9070
rect -714 9036 -678 9070
rect -644 9036 -608 9070
rect -574 9036 -538 9070
rect -504 9036 -468 9070
rect -434 9036 -398 9070
rect -364 9036 -328 9070
rect -294 9036 -258 9070
rect -224 9036 -188 9070
rect -154 9036 -118 9070
rect -84 9036 -48 9070
rect -14 9036 68 9070
rect -784 9033 68 9036
rect -784 9011 -305 9033
rect -852 9002 -305 9011
rect -271 9002 -231 9033
rect -197 9002 -157 9033
rect -123 9002 68 9033
rect -852 8939 -818 9002
rect -784 8968 -748 9002
rect -714 8968 -678 9002
rect -644 8968 -608 9002
rect -574 8968 -538 9002
rect -504 8968 -468 9002
rect -434 8968 -398 9002
rect -364 8968 -328 9002
rect -271 8999 -258 9002
rect -197 8999 -188 9002
rect -123 8999 -118 9002
rect -294 8968 -258 8999
rect -224 8968 -188 8999
rect -154 8968 -118 8999
rect -84 8968 -48 9002
rect -14 8968 68 9002
rect -784 8961 68 8968
rect -784 8939 -305 8961
rect -852 8934 -305 8939
rect -271 8934 -231 8961
rect -197 8934 -157 8961
rect -123 8934 68 8961
rect -852 8867 -818 8934
rect -784 8900 -748 8934
rect -714 8900 -678 8934
rect -644 8900 -608 8934
rect -574 8900 -538 8934
rect -504 8900 -468 8934
rect -434 8900 -398 8934
rect -364 8900 -328 8934
rect -271 8927 -258 8934
rect -197 8927 -188 8934
rect -123 8927 -118 8934
rect -294 8900 -258 8927
rect -224 8900 -188 8927
rect -154 8900 -118 8927
rect -84 8900 -48 8934
rect -14 8900 68 8934
rect -784 8889 68 8900
rect -784 8867 -305 8889
rect -852 8866 -305 8867
rect -271 8866 -231 8889
rect -197 8866 -157 8889
rect -123 8866 68 8889
rect -852 8832 -818 8866
rect -784 8832 -748 8866
rect -714 8832 -678 8866
rect -644 8832 -608 8866
rect -574 8832 -538 8866
rect -504 8832 -468 8866
rect -434 8832 -398 8866
rect -364 8832 -328 8866
rect -271 8855 -258 8866
rect -197 8855 -188 8866
rect -123 8855 -118 8866
rect -294 8832 -258 8855
rect -224 8832 -188 8855
rect -154 8832 -118 8855
rect -84 8832 -48 8866
rect -14 8832 68 8866
rect -852 8829 68 8832
rect -852 8764 -818 8829
rect -784 8817 68 8829
rect -784 8798 -305 8817
rect -271 8798 -231 8817
rect -197 8798 -157 8817
rect -123 8798 68 8817
rect -784 8764 -748 8798
rect -714 8764 -678 8798
rect -644 8764 -608 8798
rect -574 8764 -538 8798
rect -504 8764 -468 8798
rect -434 8764 -398 8798
rect -364 8764 -328 8798
rect -271 8783 -258 8798
rect -197 8783 -188 8798
rect -123 8783 -118 8798
rect -294 8764 -258 8783
rect -224 8764 -188 8783
rect -154 8764 -118 8783
rect -84 8764 -48 8798
rect -14 8764 68 8798
rect -852 8757 68 8764
rect -852 8696 -818 8757
rect -784 8745 68 8757
rect -784 8730 -305 8745
rect -271 8730 -231 8745
rect -197 8730 -157 8745
rect -123 8730 68 8745
rect -784 8696 -748 8730
rect -714 8696 -678 8730
rect -644 8696 -608 8730
rect -574 8696 -538 8730
rect -504 8696 -468 8730
rect -434 8696 -398 8730
rect -364 8696 -328 8730
rect -271 8711 -258 8730
rect -197 8711 -188 8730
rect -123 8711 -118 8730
rect -294 8696 -258 8711
rect -224 8696 -188 8711
rect -154 8696 -118 8711
rect -84 8696 -48 8730
rect -14 8696 68 8730
rect -852 8685 68 8696
rect -852 8628 -818 8685
rect -784 8673 68 8685
rect -784 8662 -305 8673
rect -271 8662 -231 8673
rect -197 8662 -157 8673
rect -123 8662 68 8673
rect -784 8628 -748 8662
rect -714 8628 -678 8662
rect -644 8628 -608 8662
rect -574 8628 -538 8662
rect -504 8628 -468 8662
rect -434 8628 -398 8662
rect -364 8628 -328 8662
rect -271 8639 -258 8662
rect -197 8639 -188 8662
rect -123 8639 -118 8662
rect -294 8628 -258 8639
rect -224 8628 -188 8639
rect -154 8628 -118 8639
rect -84 8628 -48 8662
rect -14 8628 68 8662
rect -852 8613 68 8628
rect -852 8560 -818 8613
rect -784 8601 68 8613
rect -784 8594 -305 8601
rect -271 8594 -231 8601
rect -197 8594 -157 8601
rect -123 8594 68 8601
rect -784 8560 -748 8594
rect -714 8560 -678 8594
rect -644 8560 -608 8594
rect -574 8560 -538 8594
rect -504 8560 -468 8594
rect -434 8560 -398 8594
rect -364 8560 -328 8594
rect -271 8567 -258 8594
rect -197 8567 -188 8594
rect -123 8567 -118 8594
rect -294 8560 -258 8567
rect -224 8560 -188 8567
rect -154 8560 -118 8567
rect -84 8560 -48 8594
rect -14 8560 68 8594
rect -852 8541 68 8560
rect -852 8492 -818 8541
rect -784 8529 68 8541
rect -784 8526 -305 8529
rect -271 8526 -231 8529
rect -197 8526 -157 8529
rect -123 8526 68 8529
rect -784 8492 -748 8526
rect -714 8492 -678 8526
rect -644 8492 -608 8526
rect -574 8492 -538 8526
rect -504 8492 -468 8526
rect -434 8492 -398 8526
rect -364 8492 -328 8526
rect -271 8495 -258 8526
rect -197 8495 -188 8526
rect -123 8495 -118 8526
rect -294 8492 -258 8495
rect -224 8492 -188 8495
rect -154 8492 -118 8495
rect -84 8492 -48 8526
rect -14 8492 68 8526
rect -852 8469 68 8492
rect -852 8424 -818 8469
rect -784 8458 68 8469
rect -784 8424 -748 8458
rect -714 8424 -678 8458
rect -644 8424 -608 8458
rect -574 8424 -538 8458
rect -504 8424 -468 8458
rect -434 8424 -398 8458
rect -364 8424 -328 8458
rect -294 8457 -258 8458
rect -224 8457 -188 8458
rect -154 8457 -118 8458
rect -271 8424 -258 8457
rect -197 8424 -188 8457
rect -123 8424 -118 8457
rect -84 8424 -48 8458
rect -14 8424 68 8458
rect -852 8423 -305 8424
rect -271 8423 -231 8424
rect -197 8423 -157 8424
rect -123 8423 68 8424
rect -852 8397 68 8423
rect -852 8356 -818 8397
rect -784 8390 68 8397
rect -784 8356 -748 8390
rect -714 8356 -678 8390
rect -644 8356 -608 8390
rect -574 8356 -538 8390
rect -504 8356 -468 8390
rect -434 8356 -398 8390
rect -364 8356 -328 8390
rect -294 8385 -258 8390
rect -224 8385 -188 8390
rect -154 8385 -118 8390
rect -271 8356 -258 8385
rect -197 8356 -188 8385
rect -123 8356 -118 8385
rect -84 8356 -48 8390
rect -14 8356 68 8390
rect -852 8351 -305 8356
rect -271 8351 -231 8356
rect -197 8351 -157 8356
rect -123 8351 68 8356
rect -852 8325 68 8351
rect -852 8288 -818 8325
rect -784 8322 68 8325
rect -784 8288 -748 8322
rect -714 8288 -678 8322
rect -644 8288 -608 8322
rect -574 8288 -538 8322
rect -504 8288 -468 8322
rect -434 8288 -398 8322
rect -364 8288 -328 8322
rect -294 8313 -258 8322
rect -224 8313 -188 8322
rect -154 8313 -118 8322
rect -271 8288 -258 8313
rect -197 8288 -188 8313
rect -123 8288 -118 8313
rect -84 8288 -48 8322
rect -14 8288 68 8322
rect -852 8279 -305 8288
rect -271 8279 -231 8288
rect -197 8279 -157 8288
rect -123 8279 68 8288
rect -852 8254 68 8279
rect -852 8219 -818 8254
rect -784 8220 -748 8254
rect -714 8220 -678 8254
rect -644 8220 -608 8254
rect -574 8220 -538 8254
rect -504 8220 -468 8254
rect -434 8220 -398 8254
rect -364 8220 -328 8254
rect -294 8241 -258 8254
rect -224 8241 -188 8254
rect -154 8241 -118 8254
rect -271 8220 -258 8241
rect -197 8220 -188 8241
rect -123 8220 -118 8241
rect -84 8220 -48 8254
rect -14 8220 68 8254
rect -784 8219 -305 8220
rect -852 8207 -305 8219
rect -271 8207 -231 8220
rect -197 8207 -157 8220
rect -123 8207 68 8220
rect -852 8186 68 8207
rect -852 8147 -818 8186
rect -784 8152 -748 8186
rect -714 8152 -678 8186
rect -644 8152 -608 8186
rect -574 8152 -538 8186
rect -504 8152 -468 8186
rect -434 8152 -398 8186
rect -364 8152 -328 8186
rect -294 8168 -258 8186
rect -224 8168 -188 8186
rect -154 8168 -118 8186
rect -271 8152 -258 8168
rect -197 8152 -188 8168
rect -123 8152 -118 8168
rect -84 8152 -48 8186
rect -14 8152 68 8186
rect -784 8147 -305 8152
rect -852 8134 -305 8147
rect -271 8134 -231 8152
rect -197 8134 -157 8152
rect -123 8134 68 8152
rect -852 8118 68 8134
rect -852 8075 -818 8118
rect -784 8084 -748 8118
rect -714 8084 -678 8118
rect -644 8084 -608 8118
rect -574 8084 -538 8118
rect -504 8084 -468 8118
rect -434 8084 -398 8118
rect -364 8084 -328 8118
rect -294 8095 -258 8118
rect -224 8095 -188 8118
rect -154 8095 -118 8118
rect -271 8084 -258 8095
rect -197 8084 -188 8095
rect -123 8084 -118 8095
rect -84 8084 -48 8118
rect -14 8084 68 8118
rect -784 8075 -305 8084
rect -852 8061 -305 8075
rect -271 8061 -231 8084
rect -197 8061 -157 8084
rect -123 8061 68 8084
rect -852 8050 68 8061
rect -852 8003 -818 8050
rect -784 8016 -748 8050
rect -714 8016 -678 8050
rect -644 8016 -608 8050
rect -574 8016 -538 8050
rect -504 8016 -468 8050
rect -434 8016 -398 8050
rect -364 8016 -328 8050
rect -294 8022 -258 8050
rect -224 8022 -188 8050
rect -154 8022 -118 8050
rect -271 8016 -258 8022
rect -197 8016 -188 8022
rect -123 8016 -118 8022
rect -84 8016 -48 8050
rect -14 8016 68 8050
rect -784 8003 -305 8016
rect -852 7988 -305 8003
rect -271 7988 -231 8016
rect -197 7988 -157 8016
rect -123 7988 68 8016
rect -852 7982 68 7988
rect -852 7931 -818 7982
rect -784 7948 -748 7982
rect -714 7948 -678 7982
rect -644 7948 -608 7982
rect -574 7948 -538 7982
rect -504 7948 -468 7982
rect -434 7948 -398 7982
rect -364 7948 -328 7982
rect -294 7949 -258 7982
rect -224 7949 -188 7982
rect -154 7949 -118 7982
rect -271 7948 -258 7949
rect -197 7948 -188 7949
rect -123 7948 -118 7949
rect -84 7948 -48 7982
rect -14 7948 68 7982
rect -784 7931 -305 7948
rect -852 7915 -305 7931
rect -271 7915 -231 7948
rect -197 7915 -157 7948
rect -123 7915 68 7948
rect -852 7914 68 7915
rect -852 7859 -818 7914
rect -784 7880 -748 7914
rect -714 7880 -678 7914
rect -644 7880 -608 7914
rect -574 7880 -538 7914
rect -504 7880 -468 7914
rect -434 7880 -398 7914
rect -364 7880 -328 7914
rect -294 7880 -258 7914
rect -224 7880 -188 7914
rect -154 7880 -118 7914
rect -84 7880 -48 7914
rect -14 7880 68 7914
rect -784 7876 68 7880
rect -784 7859 -305 7876
rect -852 7846 -305 7859
rect -271 7846 -231 7876
rect -197 7846 -157 7876
rect -123 7846 68 7876
rect -852 7787 -818 7846
rect -784 7812 -748 7846
rect -714 7812 -678 7846
rect -644 7812 -608 7846
rect -574 7812 -538 7846
rect -504 7812 -468 7846
rect -434 7812 -398 7846
rect -364 7812 -328 7846
rect -271 7842 -258 7846
rect -197 7842 -188 7846
rect -123 7842 -118 7846
rect -294 7812 -258 7842
rect -224 7812 -188 7842
rect -154 7812 -118 7842
rect -84 7812 -48 7846
rect -14 7812 68 7846
rect -784 7803 68 7812
rect -784 7787 -305 7803
rect -852 7778 -305 7787
rect -271 7778 -231 7803
rect -197 7778 -157 7803
rect -123 7778 68 7803
rect -852 7715 -818 7778
rect -784 7744 -748 7778
rect -714 7744 -678 7778
rect -644 7744 -608 7778
rect -574 7744 -538 7778
rect -504 7744 -468 7778
rect -434 7744 -398 7778
rect -364 7744 -328 7778
rect -271 7769 -258 7778
rect -197 7769 -188 7778
rect -123 7769 -118 7778
rect -294 7744 -258 7769
rect -224 7744 -188 7769
rect -154 7744 -118 7769
rect -84 7744 -48 7778
rect -14 7744 68 7778
rect -784 7730 68 7744
rect -784 7715 -305 7730
rect -852 7710 -305 7715
rect -271 7710 -231 7730
rect -197 7710 -157 7730
rect -123 7710 68 7730
rect -852 7643 -818 7710
rect -784 7676 -748 7710
rect -714 7676 -678 7710
rect -644 7676 -608 7710
rect -574 7676 -538 7710
rect -504 7676 -468 7710
rect -434 7676 -398 7710
rect -364 7676 -328 7710
rect -271 7696 -258 7710
rect -197 7696 -188 7710
rect -123 7696 -118 7710
rect -294 7676 -258 7696
rect -224 7676 -188 7696
rect -154 7676 -118 7696
rect -84 7676 -48 7710
rect -14 7676 68 7710
rect -784 7657 68 7676
rect -784 7643 -305 7657
rect -852 7642 -305 7643
rect -271 7642 -231 7657
rect -197 7642 -157 7657
rect -123 7642 68 7657
rect -852 7608 -818 7642
rect -784 7608 -748 7642
rect -714 7608 -678 7642
rect -644 7608 -608 7642
rect -574 7608 -538 7642
rect -504 7608 -468 7642
rect -434 7608 -398 7642
rect -364 7608 -328 7642
rect -271 7623 -258 7642
rect -197 7623 -188 7642
rect -123 7623 -118 7642
rect -294 7608 -258 7623
rect -224 7608 -188 7623
rect -154 7608 -118 7623
rect -84 7608 -48 7642
rect -14 7608 68 7642
rect -852 7605 68 7608
rect -852 7540 -818 7605
rect -784 7584 68 7605
rect -784 7574 -305 7584
rect -271 7574 -231 7584
rect -197 7574 -157 7584
rect -123 7574 68 7584
rect -784 7540 -748 7574
rect -714 7540 -678 7574
rect -644 7540 -608 7574
rect -574 7540 -538 7574
rect -504 7540 -468 7574
rect -434 7540 -398 7574
rect -364 7540 -328 7574
rect -271 7550 -258 7574
rect -197 7550 -188 7574
rect -123 7550 -118 7574
rect -294 7540 -258 7550
rect -224 7540 -188 7550
rect -154 7540 -118 7550
rect -84 7540 -48 7574
rect -14 7540 68 7574
rect -852 7533 68 7540
rect -852 7472 -818 7533
rect -784 7511 68 7533
rect -784 7506 -305 7511
rect -271 7506 -231 7511
rect -197 7506 -157 7511
rect -123 7506 68 7511
rect -784 7472 -748 7506
rect -714 7472 -678 7506
rect -644 7472 -608 7506
rect -574 7472 -538 7506
rect -504 7472 -468 7506
rect -434 7472 -398 7506
rect -364 7472 -328 7506
rect -271 7477 -258 7506
rect -197 7477 -188 7506
rect -123 7477 -118 7506
rect -294 7472 -258 7477
rect -224 7472 -188 7477
rect -154 7472 -118 7477
rect -84 7472 -48 7506
rect -14 7472 68 7506
rect -852 7461 68 7472
rect -852 7404 -818 7461
rect -784 7438 68 7461
rect -784 7404 -748 7438
rect -714 7404 -678 7438
rect -644 7404 -608 7438
rect -574 7404 -538 7438
rect -504 7404 -468 7438
rect -434 7404 -398 7438
rect -364 7404 -328 7438
rect -271 7404 -258 7438
rect -197 7404 -188 7438
rect -123 7404 -118 7438
rect -84 7404 -48 7438
rect -14 7404 68 7438
rect -852 7389 68 7404
rect -852 7336 -818 7389
rect -784 7370 68 7389
rect -784 7336 -748 7370
rect -714 7336 -678 7370
rect -644 7336 -608 7370
rect -574 7336 -538 7370
rect -504 7336 -468 7370
rect -434 7336 -398 7370
rect -364 7336 -328 7370
rect -294 7365 -258 7370
rect -224 7365 -188 7370
rect -154 7365 -118 7370
rect -271 7336 -258 7365
rect -197 7336 -188 7365
rect -123 7336 -118 7365
rect -84 7336 -48 7370
rect -14 7336 68 7370
rect -852 7331 -305 7336
rect -271 7331 -231 7336
rect -197 7331 -157 7336
rect -123 7331 68 7336
rect -852 7317 68 7331
rect -852 7268 -818 7317
rect -784 7302 68 7317
rect -784 7268 -748 7302
rect -714 7268 -678 7302
rect -644 7268 -608 7302
rect -574 7268 -538 7302
rect -504 7268 -468 7302
rect -434 7268 -398 7302
rect -364 7268 -328 7302
rect -294 7292 -258 7302
rect -224 7292 -188 7302
rect -154 7292 -118 7302
rect -271 7268 -258 7292
rect -197 7268 -188 7292
rect -123 7268 -118 7292
rect -84 7268 -48 7302
rect -14 7268 68 7302
rect -852 7258 -305 7268
rect -271 7258 -231 7268
rect -197 7258 -157 7268
rect -123 7258 68 7268
rect -852 7245 68 7258
rect -852 7200 -818 7245
rect -784 7234 68 7245
rect -784 7200 -748 7234
rect -714 7200 -678 7234
rect -644 7200 -608 7234
rect -574 7200 -538 7234
rect -504 7200 -468 7234
rect -434 7200 -398 7234
rect -364 7200 -328 7234
rect -294 7219 -258 7234
rect -224 7219 -188 7234
rect -154 7219 -118 7234
rect -271 7200 -258 7219
rect -197 7200 -188 7219
rect -123 7200 -118 7219
rect -84 7200 -48 7234
rect -14 7200 68 7234
rect -852 7185 -305 7200
rect -271 7185 -231 7200
rect -197 7185 -157 7200
rect -123 7185 68 7200
rect -852 7173 68 7185
rect -852 7132 -818 7173
rect -784 7166 68 7173
rect -784 7132 -748 7166
rect -714 7132 -678 7166
rect -644 7132 -608 7166
rect -574 7132 -538 7166
rect -504 7132 -468 7166
rect -434 7132 -398 7166
rect -364 7132 -328 7166
rect -294 7146 -258 7166
rect -224 7146 -188 7166
rect -154 7146 -118 7166
rect -271 7132 -258 7146
rect -197 7132 -188 7146
rect -123 7132 -118 7146
rect -84 7132 -48 7166
rect -14 7132 68 7166
rect -852 7112 -305 7132
rect -271 7112 -231 7132
rect -197 7112 -157 7132
rect -123 7112 68 7132
rect -852 7101 68 7112
rect -852 7064 -818 7101
rect -784 7098 68 7101
rect -784 7064 -748 7098
rect -714 7064 -678 7098
rect -644 7064 -608 7098
rect -574 7064 -538 7098
rect -504 7064 -468 7098
rect -434 7064 -398 7098
rect -364 7064 -328 7098
rect -294 7073 -258 7098
rect -224 7073 -188 7098
rect -154 7073 -118 7098
rect -271 7064 -258 7073
rect -197 7064 -188 7073
rect -123 7064 -118 7073
rect -84 7064 -48 7098
rect -14 7064 68 7098
rect -852 7039 -305 7064
rect -271 7039 -231 7064
rect -197 7039 -157 7064
rect -123 7039 68 7064
rect -852 7030 68 7039
rect -852 6995 -818 7030
rect -784 6996 -748 7030
rect -714 6996 -678 7030
rect -644 6996 -608 7030
rect -574 6996 -538 7030
rect -504 6996 -468 7030
rect -434 6996 -398 7030
rect -364 6996 -328 7030
rect -294 7000 -258 7030
rect -224 7000 -188 7030
rect -154 7000 -118 7030
rect -271 6996 -258 7000
rect -197 6996 -188 7000
rect -123 6996 -118 7000
rect -84 6996 -48 7030
rect -14 6996 68 7030
rect -784 6995 -305 6996
rect -852 6966 -305 6995
rect -271 6966 -231 6996
rect -197 6966 -157 6996
rect -123 6966 68 6996
rect -852 6962 68 6966
rect -852 6923 -818 6962
rect -784 6928 -748 6962
rect -714 6928 -678 6962
rect -644 6928 -608 6962
rect -574 6928 -538 6962
rect -504 6928 -468 6962
rect -434 6928 -398 6962
rect -364 6928 -328 6962
rect -294 6928 -258 6962
rect -224 6928 -188 6962
rect -154 6928 -118 6962
rect -84 6928 -48 6962
rect -14 6928 68 6962
rect -784 6927 68 6928
rect -784 6923 -305 6927
rect -852 6894 -305 6923
rect -271 6894 -231 6927
rect -197 6894 -157 6927
rect -123 6894 68 6927
rect -852 6851 -818 6894
rect -784 6860 -748 6894
rect -714 6860 -678 6894
rect -644 6860 -608 6894
rect -574 6860 -538 6894
rect -504 6860 -468 6894
rect -434 6860 -398 6894
rect -364 6860 -328 6894
rect -271 6893 -258 6894
rect -197 6893 -188 6894
rect -123 6893 -118 6894
rect -294 6860 -258 6893
rect -224 6860 -188 6893
rect -154 6860 -118 6893
rect -84 6860 -48 6894
rect -14 6860 68 6894
rect -784 6854 68 6860
rect -784 6851 -305 6854
rect -852 6826 -305 6851
rect -271 6826 -231 6854
rect -197 6826 -157 6854
rect -123 6826 68 6854
rect -852 6779 -818 6826
rect -784 6792 -748 6826
rect -714 6792 -678 6826
rect -644 6792 -608 6826
rect -574 6792 -538 6826
rect -504 6792 -468 6826
rect -434 6792 -398 6826
rect -364 6792 -328 6826
rect -271 6820 -258 6826
rect -197 6820 -188 6826
rect -123 6820 -118 6826
rect -294 6792 -258 6820
rect -224 6792 -188 6820
rect -154 6792 -118 6820
rect -84 6792 -48 6826
rect -14 6792 68 6826
rect -784 6781 68 6792
rect -784 6779 -305 6781
rect -852 6758 -305 6779
rect -271 6758 -231 6781
rect -197 6758 -157 6781
rect -123 6758 68 6781
rect -852 6707 -818 6758
rect -784 6724 -748 6758
rect -714 6724 -678 6758
rect -644 6724 -608 6758
rect -574 6724 -538 6758
rect -504 6724 -468 6758
rect -434 6724 -398 6758
rect -364 6724 -328 6758
rect -271 6747 -258 6758
rect -197 6747 -188 6758
rect -123 6747 -118 6758
rect -294 6724 -258 6747
rect -224 6724 -188 6747
rect -154 6724 -118 6747
rect -84 6724 -48 6758
rect -14 6724 68 6758
rect -784 6708 68 6724
rect -784 6707 -305 6708
rect -852 6690 -305 6707
rect -271 6690 -231 6708
rect -197 6690 -157 6708
rect -123 6690 68 6708
rect -852 6635 -818 6690
rect -784 6656 -748 6690
rect -714 6656 -678 6690
rect -644 6656 -608 6690
rect -574 6656 -538 6690
rect -504 6656 -468 6690
rect -434 6656 -398 6690
rect -364 6656 -328 6690
rect -271 6674 -258 6690
rect -197 6674 -188 6690
rect -123 6674 -118 6690
rect -294 6656 -258 6674
rect -224 6656 -188 6674
rect -154 6656 -118 6674
rect -84 6656 -48 6690
rect -14 6656 68 6690
rect -784 6635 68 6656
rect -852 6622 -305 6635
rect -271 6622 -231 6635
rect -197 6622 -157 6635
rect -123 6622 68 6635
rect -852 6563 -818 6622
rect -784 6588 -748 6622
rect -714 6588 -678 6622
rect -644 6588 -608 6622
rect -574 6588 -538 6622
rect -504 6588 -468 6622
rect -434 6588 -398 6622
rect -364 6588 -328 6622
rect -271 6601 -258 6622
rect -197 6601 -188 6622
rect -123 6601 -118 6622
rect -294 6588 -258 6601
rect -224 6588 -188 6601
rect -154 6588 -118 6601
rect -84 6588 -48 6622
rect -14 6588 68 6622
rect -784 6563 68 6588
rect -852 6562 68 6563
rect -852 6554 -305 6562
rect -271 6554 -231 6562
rect -197 6554 -157 6562
rect -123 6554 68 6562
rect -852 6491 -818 6554
rect -784 6520 -748 6554
rect -714 6520 -678 6554
rect -644 6520 -608 6554
rect -574 6520 -538 6554
rect -504 6520 -468 6554
rect -434 6520 -398 6554
rect -364 6520 -328 6554
rect -271 6528 -258 6554
rect -197 6528 -188 6554
rect -123 6528 -118 6554
rect -294 6520 -258 6528
rect -224 6520 -188 6528
rect -154 6520 -118 6528
rect -84 6520 -48 6554
rect -14 6520 68 6554
rect -784 6491 68 6520
rect -852 6489 68 6491
rect -852 6486 -305 6489
rect -271 6486 -231 6489
rect -197 6486 -157 6489
rect -123 6486 68 6489
rect -852 6419 -818 6486
rect -784 6452 -748 6486
rect -714 6452 -678 6486
rect -644 6452 -608 6486
rect -574 6452 -538 6486
rect -504 6452 -468 6486
rect -434 6452 -398 6486
rect -364 6452 -328 6486
rect -271 6455 -258 6486
rect -197 6455 -188 6486
rect -123 6455 -118 6486
rect -294 6452 -258 6455
rect -224 6452 -188 6455
rect -154 6452 -118 6455
rect -84 6452 -48 6486
rect -14 6452 68 6486
rect -784 6419 68 6452
rect -852 6418 68 6419
rect -852 6384 -818 6418
rect -784 6384 -748 6418
rect -714 6384 -678 6418
rect -644 6384 -608 6418
rect -574 6384 -538 6418
rect -504 6384 -468 6418
rect -434 6384 -398 6418
rect -364 6384 -328 6418
rect -294 6416 -258 6418
rect -224 6416 -188 6418
rect -154 6416 -118 6418
rect -271 6384 -258 6416
rect -197 6384 -188 6416
rect -123 6384 -118 6416
rect -84 6384 -48 6418
rect -14 6384 68 6418
rect -852 6382 -305 6384
rect -271 6382 -231 6384
rect -197 6382 -157 6384
rect -123 6382 68 6384
rect -852 6381 68 6382
rect -852 6316 -818 6381
rect -784 6350 68 6381
rect -784 6316 -748 6350
rect -714 6316 -678 6350
rect -644 6316 -608 6350
rect -574 6316 -538 6350
rect -504 6316 -468 6350
rect -434 6316 -398 6350
rect -364 6316 -328 6350
rect -294 6343 -258 6350
rect -224 6343 -188 6350
rect -154 6343 -118 6350
rect -271 6316 -258 6343
rect -197 6316 -188 6343
rect -123 6316 -118 6343
rect -84 6316 -48 6350
rect -14 6316 68 6350
rect -852 6309 -305 6316
rect -271 6309 -231 6316
rect -197 6309 -157 6316
rect -123 6309 68 6316
rect -852 6248 -818 6309
rect -784 6282 68 6309
rect -784 6248 -748 6282
rect -714 6248 -678 6282
rect -644 6248 -608 6282
rect -574 6248 -538 6282
rect -504 6248 -468 6282
rect -434 6248 -398 6282
rect -364 6248 -328 6282
rect -294 6270 -258 6282
rect -224 6270 -188 6282
rect -154 6270 -118 6282
rect -271 6248 -258 6270
rect -197 6248 -188 6270
rect -123 6248 -118 6270
rect -84 6248 -48 6282
rect -14 6248 68 6282
rect -852 6237 -305 6248
rect -852 6180 -818 6237
rect -784 6236 -305 6237
rect -271 6236 -231 6248
rect -197 6236 -157 6248
rect -123 6236 68 6248
rect -784 6214 68 6236
rect -784 6180 -748 6214
rect -714 6180 -678 6214
rect -644 6180 -608 6214
rect -574 6180 -538 6214
rect -504 6180 -468 6214
rect -434 6180 -398 6214
rect -364 6180 -328 6214
rect -294 6197 -258 6214
rect -224 6197 -188 6214
rect -154 6197 -118 6214
rect -271 6180 -258 6197
rect -197 6180 -188 6197
rect -123 6180 -118 6197
rect -84 6180 -48 6214
rect -14 6180 68 6214
rect -852 6165 -305 6180
rect -852 6112 -818 6165
rect -784 6163 -305 6165
rect -271 6163 -231 6180
rect -197 6163 -157 6180
rect -123 6163 68 6180
rect -784 6146 68 6163
rect -784 6112 -748 6146
rect -714 6112 -678 6146
rect -644 6112 -608 6146
rect -574 6112 -538 6146
rect -504 6112 -468 6146
rect -434 6112 -398 6146
rect -364 6112 -328 6146
rect -294 6124 -258 6146
rect -224 6124 -188 6146
rect -154 6124 -118 6146
rect -271 6112 -258 6124
rect -197 6112 -188 6124
rect -123 6112 -118 6124
rect -84 6112 -48 6146
rect -14 6112 68 6146
rect -852 6093 -305 6112
rect -852 6044 -818 6093
rect -784 6090 -305 6093
rect -271 6090 -231 6112
rect -197 6090 -157 6112
rect -123 6090 68 6112
rect -784 6078 68 6090
rect -784 6044 -748 6078
rect -714 6044 -678 6078
rect -644 6044 -608 6078
rect -574 6044 -538 6078
rect -504 6044 -468 6078
rect -434 6044 -398 6078
rect -364 6044 -328 6078
rect -294 6051 -258 6078
rect -224 6051 -188 6078
rect -154 6051 -118 6078
rect -271 6044 -258 6051
rect -197 6044 -188 6051
rect -123 6044 -118 6051
rect -84 6044 -48 6078
rect -14 6044 68 6078
rect -852 6021 -305 6044
rect -852 5976 -818 6021
rect -784 6017 -305 6021
rect -271 6017 -231 6044
rect -197 6017 -157 6044
rect -123 6017 68 6044
rect -784 6010 68 6017
rect -784 5976 -748 6010
rect -714 5976 -678 6010
rect -644 5976 -608 6010
rect -574 5976 -538 6010
rect -504 5976 -468 6010
rect -434 5976 -398 6010
rect -364 5976 -328 6010
rect -294 5978 -258 6010
rect -224 5978 -188 6010
rect -154 5978 -118 6010
rect -271 5976 -258 5978
rect -197 5976 -188 5978
rect -123 5976 -118 5978
rect -84 5976 -48 6010
rect -14 5976 68 6010
rect -852 5949 -305 5976
rect -852 5908 -818 5949
rect -784 5944 -305 5949
rect -271 5944 -231 5976
rect -197 5944 -157 5976
rect -123 5944 68 5976
rect -784 5942 68 5944
rect -784 5908 -748 5942
rect -714 5908 -678 5942
rect -644 5908 -608 5942
rect -574 5908 -538 5942
rect -504 5908 -468 5942
rect -434 5908 -398 5942
rect -364 5908 -328 5942
rect -294 5908 -258 5942
rect -224 5908 -188 5942
rect -154 5908 -118 5942
rect -84 5908 -48 5942
rect -14 5908 68 5942
rect -852 5905 68 5908
rect -852 5877 -305 5905
rect -852 5840 -818 5877
rect -784 5874 -305 5877
rect -271 5874 -231 5905
rect -197 5874 -157 5905
rect -123 5874 68 5905
rect -784 5840 -748 5874
rect -714 5840 -678 5874
rect -644 5840 -608 5874
rect -574 5840 -538 5874
rect -504 5840 -468 5874
rect -434 5840 -398 5874
rect -364 5840 -328 5874
rect -271 5871 -258 5874
rect -197 5871 -188 5874
rect -123 5871 -118 5874
rect -294 5840 -258 5871
rect -224 5840 -188 5871
rect -154 5840 -118 5871
rect -84 5840 -48 5874
rect -14 5840 68 5874
rect -852 5832 68 5840
rect -852 5806 -305 5832
rect -271 5806 -231 5832
rect -197 5806 -157 5832
rect -123 5806 68 5832
rect -852 5771 -818 5806
rect -784 5772 -748 5806
rect -714 5772 -678 5806
rect -644 5772 -608 5806
rect -574 5772 -538 5806
rect -504 5772 -468 5806
rect -434 5772 -398 5806
rect -364 5772 -328 5806
rect -271 5798 -258 5806
rect -197 5798 -188 5806
rect -123 5798 -118 5806
rect -294 5772 -258 5798
rect -224 5772 -188 5798
rect -154 5772 -118 5798
rect -84 5772 -48 5806
rect -14 5772 68 5806
rect -784 5771 68 5772
rect -852 5759 68 5771
rect -852 5738 -305 5759
rect -271 5738 -231 5759
rect -197 5738 -157 5759
rect -123 5738 68 5759
rect -852 5699 -818 5738
rect -784 5704 -748 5738
rect -714 5704 -678 5738
rect -644 5704 -608 5738
rect -574 5704 -538 5738
rect -504 5704 -468 5738
rect -434 5704 -398 5738
rect -364 5704 -328 5738
rect -271 5725 -258 5738
rect -197 5725 -188 5738
rect -123 5725 -118 5738
rect -294 5704 -258 5725
rect -224 5704 -188 5725
rect -154 5704 -118 5725
rect -84 5704 -48 5738
rect -14 5704 68 5738
rect -784 5699 68 5704
rect -852 5686 68 5699
rect -852 5670 -305 5686
rect -271 5670 -231 5686
rect -197 5670 -157 5686
rect -123 5670 68 5686
rect -852 5627 -818 5670
rect -784 5636 -748 5670
rect -714 5636 -678 5670
rect -644 5636 -608 5670
rect -574 5636 -538 5670
rect -504 5636 -468 5670
rect -434 5636 -398 5670
rect -364 5636 -328 5670
rect -271 5652 -258 5670
rect -197 5652 -188 5670
rect -123 5652 -118 5670
rect -294 5636 -258 5652
rect -224 5636 -188 5652
rect -154 5636 -118 5652
rect -84 5636 -48 5670
rect -14 5636 68 5670
rect -784 5627 68 5636
rect -852 5613 68 5627
rect -852 5602 -305 5613
rect -271 5602 -231 5613
rect -197 5602 -157 5613
rect -123 5602 68 5613
rect -852 5555 -818 5602
rect -784 5568 -748 5602
rect -714 5568 -678 5602
rect -644 5568 -608 5602
rect -574 5568 -538 5602
rect -504 5568 -468 5602
rect -434 5568 -398 5602
rect -364 5568 -328 5602
rect -271 5579 -258 5602
rect -197 5579 -188 5602
rect -123 5579 -118 5602
rect -294 5568 -258 5579
rect -224 5568 -188 5579
rect -154 5568 -118 5579
rect -84 5568 -48 5602
rect -14 5568 68 5602
rect -784 5555 68 5568
rect -852 5540 68 5555
rect -852 5534 -305 5540
rect -271 5534 -231 5540
rect -197 5534 -157 5540
rect -123 5534 68 5540
rect -852 5483 -818 5534
rect -784 5500 -748 5534
rect -714 5500 -678 5534
rect -644 5500 -608 5534
rect -574 5500 -538 5534
rect -504 5500 -468 5534
rect -434 5500 -398 5534
rect -364 5500 -328 5534
rect -271 5506 -258 5534
rect -197 5506 -188 5534
rect -123 5506 -118 5534
rect -294 5500 -258 5506
rect -224 5500 -188 5506
rect -154 5500 -118 5506
rect -84 5500 -48 5534
rect -14 5500 68 5534
rect -784 5483 68 5500
rect -852 5467 68 5483
rect -852 5466 -305 5467
rect -271 5466 -231 5467
rect -197 5466 -157 5467
rect -123 5466 68 5467
rect -852 5411 -818 5466
rect -784 5432 -748 5466
rect -714 5432 -678 5466
rect -644 5432 -608 5466
rect -574 5432 -538 5466
rect -504 5432 -468 5466
rect -434 5432 -398 5466
rect -364 5432 -328 5466
rect -271 5433 -258 5466
rect -197 5433 -188 5466
rect -123 5433 -118 5466
rect -294 5432 -258 5433
rect -224 5432 -188 5433
rect -154 5432 -118 5433
rect -84 5432 -48 5466
rect -14 5432 68 5466
rect -784 5411 68 5432
rect -852 5398 68 5411
rect -852 5339 -818 5398
rect -784 5364 -748 5398
rect -714 5364 -678 5398
rect -644 5364 -608 5398
rect -574 5364 -538 5398
rect -504 5364 -468 5398
rect -434 5364 -398 5398
rect -364 5364 -328 5398
rect -294 5394 -258 5398
rect -224 5394 -188 5398
rect -154 5394 -118 5398
rect -271 5364 -258 5394
rect -197 5364 -188 5394
rect -123 5364 -118 5394
rect -84 5364 -48 5398
rect -14 5364 68 5398
rect -784 5360 -305 5364
rect -271 5360 -231 5364
rect -197 5360 -157 5364
rect -123 5360 68 5364
rect -784 5339 68 5360
rect -852 5330 68 5339
rect -852 5267 -818 5330
rect -784 5296 -748 5330
rect -714 5296 -678 5330
rect -644 5296 -608 5330
rect -574 5296 -538 5330
rect -504 5296 -468 5330
rect -434 5296 -398 5330
rect -364 5296 -328 5330
rect -294 5321 -258 5330
rect -224 5321 -188 5330
rect -154 5321 -118 5330
rect -271 5296 -258 5321
rect -197 5296 -188 5321
rect -123 5296 -118 5321
rect -84 5296 -48 5330
rect -14 5296 68 5330
rect -784 5287 -305 5296
rect -271 5287 -231 5296
rect -197 5287 -157 5296
rect -123 5287 68 5296
rect -784 5267 68 5287
rect -852 5262 68 5267
rect -852 5195 -818 5262
rect -784 5228 -748 5262
rect -714 5228 -678 5262
rect -644 5228 -608 5262
rect -574 5228 -538 5262
rect -504 5228 -468 5262
rect -434 5228 -398 5262
rect -364 5228 -328 5262
rect -294 5248 -258 5262
rect -224 5248 -188 5262
rect -154 5248 -118 5262
rect -271 5228 -258 5248
rect -197 5228 -188 5248
rect -123 5228 -118 5248
rect -84 5228 -48 5262
rect -14 5228 68 5262
rect -784 5214 -305 5228
rect -271 5214 -231 5228
rect -197 5214 -157 5228
rect -123 5214 68 5228
rect -784 5195 68 5214
rect -852 5194 68 5195
rect -852 5160 -818 5194
rect -784 5160 -748 5194
rect -714 5160 -678 5194
rect -644 5160 -608 5194
rect -574 5160 -538 5194
rect -504 5160 -468 5194
rect -434 5160 -398 5194
rect -364 5160 -328 5194
rect -294 5175 -258 5194
rect -224 5175 -188 5194
rect -154 5175 -118 5194
rect -271 5160 -258 5175
rect -197 5160 -188 5175
rect -123 5160 -118 5175
rect -84 5160 -48 5194
rect -14 5160 68 5194
rect -852 5157 -305 5160
rect -852 5092 -818 5157
rect -784 5141 -305 5157
rect -271 5141 -231 5160
rect -197 5141 -157 5160
rect -123 5141 68 5160
rect -784 5126 68 5141
rect -784 5092 -748 5126
rect -714 5092 -678 5126
rect -644 5092 -608 5126
rect -574 5092 -538 5126
rect -504 5092 -468 5126
rect -434 5092 -398 5126
rect -364 5092 -328 5126
rect -294 5102 -258 5126
rect -224 5102 -188 5126
rect -154 5102 -118 5126
rect -271 5092 -258 5102
rect -197 5092 -188 5102
rect -123 5092 -118 5102
rect -84 5092 -48 5126
rect -14 5092 68 5126
rect -852 5085 -305 5092
rect -852 5024 -818 5085
rect -784 5068 -305 5085
rect -271 5068 -231 5092
rect -197 5068 -157 5092
rect -123 5068 68 5092
rect -784 5058 68 5068
rect -784 5024 -748 5058
rect -714 5024 -678 5058
rect -644 5024 -608 5058
rect -574 5024 -538 5058
rect -504 5024 -468 5058
rect -434 5024 -398 5058
rect -364 5024 -328 5058
rect -294 5029 -258 5058
rect -224 5029 -188 5058
rect -154 5029 -118 5058
rect -271 5024 -258 5029
rect -197 5024 -188 5029
rect -123 5024 -118 5029
rect -84 5024 -48 5058
rect -14 5024 68 5058
rect -852 5013 -305 5024
rect -852 4956 -818 5013
rect -784 4995 -305 5013
rect -271 4995 -231 5024
rect -197 4995 -157 5024
rect -123 5010 68 5024
rect -123 4995 28 5010
rect -784 4990 28 4995
rect -784 4956 -748 4990
rect -714 4956 -678 4990
rect -644 4956 -608 4990
rect -574 4956 -538 4990
rect -504 4956 -468 4990
rect -434 4956 -398 4990
rect -364 4956 -328 4990
rect -294 4956 -258 4990
rect -224 4956 -188 4990
rect -154 4956 -118 4990
rect -84 4974 -48 4990
rect -14 4976 28 4990
rect 62 4986 106 5010
rect 62 4976 68 4986
rect -84 4956 -62 4974
rect -14 4956 68 4976
rect -852 4941 -305 4956
rect -852 4888 -818 4941
rect -784 4922 -305 4941
rect -271 4922 -231 4956
rect -197 4922 -157 4956
rect -123 4940 -62 4956
rect -28 4952 68 4956
rect 102 4976 106 4986
rect 140 4976 184 5010
rect 218 4976 262 5010
rect 296 4976 340 5010
rect 374 4976 418 5010
rect 452 4976 496 5010
rect 530 4976 574 5010
rect 608 4976 652 5010
rect 686 4976 730 5010
rect 764 4976 808 5010
rect 842 4976 882 5010
rect -28 4940 102 4952
rect -123 4922 102 4940
rect -784 4888 -748 4922
rect -714 4888 -678 4922
rect -644 4888 -608 4922
rect -574 4888 -538 4922
rect -504 4888 -468 4922
rect -434 4888 -398 4922
rect -364 4888 -328 4922
rect -294 4888 -258 4922
rect -224 4888 -188 4922
rect -154 4888 -118 4922
rect -84 4901 -48 4922
rect -14 4918 102 4922
rect -84 4888 -62 4901
rect -14 4888 68 4918
rect -852 4883 -62 4888
rect -852 4869 -305 4883
rect -852 4820 -818 4869
rect -784 4854 -305 4869
rect -271 4854 -231 4883
rect -197 4854 -157 4883
rect -123 4867 -62 4883
rect -28 4884 68 4888
rect -28 4867 102 4884
rect -123 4854 102 4867
rect -784 4820 -748 4854
rect -714 4820 -678 4854
rect -644 4820 -608 4854
rect -574 4820 -538 4854
rect -504 4820 -468 4854
rect -434 4820 -398 4854
rect -364 4820 -328 4854
rect -271 4849 -258 4854
rect -197 4849 -188 4854
rect -123 4849 -118 4854
rect -294 4820 -258 4849
rect -224 4820 -188 4849
rect -154 4820 -118 4849
rect -84 4828 -48 4854
rect -14 4850 102 4854
rect -84 4820 -62 4828
rect -14 4820 68 4850
rect -852 4810 -62 4820
rect -852 4797 -305 4810
rect -852 4752 -818 4797
rect -784 4786 -305 4797
rect -271 4786 -231 4810
rect -197 4786 -157 4810
rect -123 4794 -62 4810
rect -28 4816 68 4820
rect -28 4794 102 4816
rect -123 4786 102 4794
rect -784 4752 -748 4786
rect -714 4752 -678 4786
rect -644 4752 -608 4786
rect -574 4752 -538 4786
rect -504 4752 -468 4786
rect -434 4752 -398 4786
rect -364 4752 -328 4786
rect -271 4776 -258 4786
rect -197 4776 -188 4786
rect -123 4776 -118 4786
rect -294 4752 -258 4776
rect -224 4752 -188 4776
rect -154 4752 -118 4776
rect -84 4755 -48 4786
rect -14 4782 102 4786
rect -84 4752 -62 4755
rect -14 4752 68 4782
rect -852 4737 -62 4752
rect -852 4725 -305 4737
rect -852 4684 -818 4725
rect -784 4718 -305 4725
rect -271 4718 -231 4737
rect -197 4718 -157 4737
rect -123 4721 -62 4737
rect -28 4748 68 4752
rect -28 4721 102 4748
rect -123 4718 102 4721
rect -784 4684 -748 4718
rect -714 4684 -678 4718
rect -644 4684 -608 4718
rect -574 4684 -538 4718
rect -504 4684 -468 4718
rect -434 4684 -398 4718
rect -364 4684 -328 4718
rect -271 4703 -258 4718
rect -197 4703 -188 4718
rect -123 4703 -118 4718
rect -294 4684 -258 4703
rect -224 4684 -188 4703
rect -154 4684 -118 4703
rect -84 4684 -48 4718
rect -14 4714 102 4718
rect -14 4684 68 4714
rect -852 4682 68 4684
rect -852 4664 -62 4682
rect -852 4653 -305 4664
rect -852 4616 -818 4653
rect -784 4650 -305 4653
rect -271 4650 -231 4664
rect -197 4650 -157 4664
rect -123 4650 -62 4664
rect -28 4680 68 4682
rect -28 4650 102 4680
rect -784 4616 -748 4650
rect -714 4616 -678 4650
rect -644 4616 -608 4650
rect -574 4616 -538 4650
rect -504 4616 -468 4650
rect -434 4616 -398 4650
rect -364 4616 -328 4650
rect -271 4630 -258 4650
rect -197 4630 -188 4650
rect -123 4630 -118 4650
rect -294 4616 -258 4630
rect -224 4616 -188 4630
rect -154 4616 -118 4630
rect -84 4648 -62 4650
rect -84 4616 -48 4648
rect -14 4646 102 4650
rect -14 4616 68 4646
rect -852 4612 68 4616
rect -852 4609 102 4612
rect -852 4591 -62 4609
rect -852 4582 -305 4591
rect -271 4582 -231 4591
rect -197 4582 -157 4591
rect -123 4582 -62 4591
rect -28 4582 102 4609
rect -852 4547 -818 4582
rect -784 4548 -748 4582
rect -714 4548 -678 4582
rect -644 4548 -608 4582
rect -574 4548 -538 4582
rect -504 4548 -468 4582
rect -434 4548 -398 4582
rect -364 4548 -328 4582
rect -271 4557 -258 4582
rect -197 4557 -188 4582
rect -123 4557 -118 4582
rect -294 4548 -258 4557
rect -224 4548 -188 4557
rect -154 4548 -118 4557
rect -84 4575 -62 4582
rect -14 4578 102 4582
rect -84 4548 -48 4575
rect -14 4548 68 4578
rect -784 4547 68 4548
rect -852 4544 68 4547
rect -852 4536 102 4544
rect -852 4518 -62 4536
rect -852 4514 -305 4518
rect -271 4514 -231 4518
rect -197 4514 -157 4518
rect -123 4514 -62 4518
rect -28 4514 102 4536
rect -852 4475 -818 4514
rect -784 4480 -748 4514
rect -714 4480 -678 4514
rect -644 4480 -608 4514
rect -574 4480 -538 4514
rect -504 4480 -468 4514
rect -434 4480 -398 4514
rect -364 4480 -328 4514
rect -271 4484 -258 4514
rect -197 4484 -188 4514
rect -123 4484 -118 4514
rect -294 4480 -258 4484
rect -224 4480 -188 4484
rect -154 4480 -118 4484
rect -84 4502 -62 4514
rect -14 4510 102 4514
rect -84 4480 -48 4502
rect -14 4480 68 4510
rect -784 4476 68 4480
rect -784 4475 102 4476
rect -852 4463 102 4475
rect -852 4446 -62 4463
rect -28 4446 102 4463
rect -852 4403 -818 4446
rect -784 4412 -748 4446
rect -714 4412 -678 4446
rect -644 4412 -608 4446
rect -574 4412 -538 4446
rect -504 4412 -468 4446
rect -434 4412 -398 4446
rect -364 4412 -328 4446
rect -294 4445 -258 4446
rect -224 4445 -188 4446
rect -154 4445 -118 4446
rect -271 4412 -258 4445
rect -197 4412 -188 4445
rect -123 4412 -118 4445
rect -84 4429 -62 4446
rect -14 4442 102 4446
rect -84 4412 -48 4429
rect -14 4412 68 4442
rect -784 4411 -305 4412
rect -271 4411 -231 4412
rect -197 4411 -157 4412
rect -123 4411 68 4412
rect -784 4408 68 4411
rect -784 4403 102 4408
rect -852 4390 102 4403
rect -852 4378 -62 4390
rect -28 4378 102 4390
rect -852 4331 -818 4378
rect -784 4344 -748 4378
rect -714 4344 -678 4378
rect -644 4344 -608 4378
rect -574 4344 -538 4378
rect -504 4344 -468 4378
rect -434 4344 -398 4378
rect -364 4344 -328 4378
rect -294 4372 -258 4378
rect -224 4372 -188 4378
rect -154 4372 -118 4378
rect -271 4344 -258 4372
rect -197 4344 -188 4372
rect -123 4344 -118 4372
rect -84 4356 -62 4378
rect -14 4374 102 4378
rect -84 4344 -48 4356
rect -14 4344 68 4374
rect -784 4338 -305 4344
rect -271 4338 -231 4344
rect -197 4338 -157 4344
rect -123 4340 68 4344
rect -123 4338 102 4340
rect -784 4331 102 4338
rect -852 4317 102 4331
rect -852 4310 -62 4317
rect -28 4310 102 4317
rect -852 4259 -818 4310
rect -784 4276 -748 4310
rect -714 4276 -678 4310
rect -644 4276 -608 4310
rect -574 4276 -538 4310
rect -504 4276 -468 4310
rect -434 4276 -398 4310
rect -364 4276 -328 4310
rect -294 4299 -258 4310
rect -224 4299 -188 4310
rect -154 4299 -118 4310
rect -271 4276 -258 4299
rect -197 4276 -188 4299
rect -123 4276 -118 4299
rect -84 4283 -62 4310
rect -14 4306 102 4310
rect -84 4276 -48 4283
rect -14 4276 68 4306
rect -784 4265 -305 4276
rect -271 4265 -231 4276
rect -197 4265 -157 4276
rect -123 4272 68 4276
rect -123 4265 102 4272
rect -784 4259 102 4265
rect -852 4244 102 4259
rect -852 4242 -62 4244
rect -28 4242 102 4244
rect -852 4187 -818 4242
rect -784 4208 -748 4242
rect -714 4208 -678 4242
rect -644 4208 -608 4242
rect -574 4208 -538 4242
rect -504 4208 -468 4242
rect -434 4208 -398 4242
rect -364 4208 -328 4242
rect -294 4226 -258 4242
rect -224 4226 -188 4242
rect -154 4226 -118 4242
rect -271 4208 -258 4226
rect -197 4208 -188 4226
rect -123 4208 -118 4226
rect -84 4210 -62 4242
rect -14 4238 102 4242
rect -84 4208 -48 4210
rect -14 4208 68 4238
rect -784 4192 -305 4208
rect -271 4192 -231 4208
rect -197 4192 -157 4208
rect -123 4204 68 4208
rect -123 4192 102 4204
rect -784 4187 102 4192
rect -852 4174 102 4187
rect -852 4115 -818 4174
rect -784 4140 -748 4174
rect -714 4140 -678 4174
rect -644 4140 -608 4174
rect -574 4140 -538 4174
rect -504 4140 -468 4174
rect -434 4140 -398 4174
rect -364 4140 -328 4174
rect -294 4153 -258 4174
rect -224 4153 -188 4174
rect -154 4153 -118 4174
rect -271 4140 -258 4153
rect -197 4140 -188 4153
rect -123 4140 -118 4153
rect -84 4171 -48 4174
rect -84 4140 -62 4171
rect -14 4170 102 4174
rect -14 4140 68 4170
rect -784 4119 -305 4140
rect -271 4119 -231 4140
rect -197 4119 -157 4140
rect -123 4137 -62 4140
rect -28 4137 68 4140
rect -123 4136 68 4137
rect -123 4119 102 4136
rect -784 4115 102 4119
rect -852 4106 102 4115
rect -852 4043 -818 4106
rect -784 4072 -748 4106
rect -714 4072 -678 4106
rect -644 4072 -608 4106
rect -574 4072 -538 4106
rect -504 4072 -468 4106
rect -434 4072 -398 4106
rect -364 4072 -328 4106
rect -294 4080 -258 4106
rect -224 4080 -188 4106
rect -154 4080 -118 4106
rect -271 4072 -258 4080
rect -197 4072 -188 4080
rect -123 4072 -118 4080
rect -84 4098 -48 4106
rect -14 4102 102 4106
rect -84 4072 -62 4098
rect -14 4072 68 4102
rect -784 4046 -305 4072
rect -271 4046 -231 4072
rect -197 4046 -157 4072
rect -123 4064 -62 4072
rect -28 4068 68 4072
rect -28 4064 102 4068
rect -123 4046 102 4064
rect -784 4043 102 4046
rect -852 4038 102 4043
rect -852 3971 -818 4038
rect -784 4004 -748 4038
rect -714 4004 -678 4038
rect -644 4004 -608 4038
rect -574 4004 -538 4038
rect -504 4004 -468 4038
rect -434 4004 -398 4038
rect -364 4004 -328 4038
rect -294 4007 -258 4038
rect -224 4007 -188 4038
rect -154 4007 -118 4038
rect -271 4004 -258 4007
rect -197 4004 -188 4007
rect -123 4004 -118 4007
rect -84 4026 -48 4038
rect -14 4034 102 4038
rect -84 4004 -62 4026
rect -14 4004 68 4034
rect -784 3973 -305 4004
rect -271 3973 -231 4004
rect -197 3973 -157 4004
rect -123 3992 -62 4004
rect -28 4000 68 4004
rect -28 3992 102 4000
rect -123 3973 102 3992
rect -784 3971 102 3973
rect -852 3970 102 3971
rect -852 3936 -818 3970
rect -784 3936 -748 3970
rect -714 3936 -678 3970
rect -644 3936 -608 3970
rect -574 3936 -538 3970
rect -504 3936 -468 3970
rect -434 3936 -398 3970
rect -364 3936 -328 3970
rect -294 3936 -258 3970
rect -224 3936 -188 3970
rect -154 3936 -118 3970
rect -84 3954 -48 3970
rect -14 3966 102 3970
rect -84 3936 -62 3954
rect -14 3936 68 3966
rect -852 3934 -62 3936
rect -852 3933 -305 3934
rect -852 3868 -818 3933
rect -784 3902 -305 3933
rect -271 3902 -231 3934
rect -197 3902 -157 3934
rect -123 3920 -62 3934
rect -28 3932 68 3936
rect -28 3920 102 3932
rect -123 3902 102 3920
rect -784 3868 -748 3902
rect -714 3868 -678 3902
rect -644 3868 -608 3902
rect -574 3868 -538 3902
rect -504 3868 -468 3902
rect -434 3868 -398 3902
rect -364 3868 -328 3902
rect -271 3900 -258 3902
rect -197 3900 -188 3902
rect -123 3900 -118 3902
rect -294 3868 -258 3900
rect -224 3868 -188 3900
rect -154 3868 -118 3900
rect -84 3882 -48 3902
rect -14 3898 102 3902
rect -84 3868 -62 3882
rect -14 3868 68 3898
rect -852 3861 -62 3868
rect -852 3800 -818 3861
rect -784 3834 -305 3861
rect -271 3834 -231 3861
rect -197 3834 -157 3861
rect -123 3848 -62 3861
rect -28 3864 68 3868
rect -28 3848 102 3864
rect -123 3834 102 3848
rect -784 3800 -748 3834
rect -714 3800 -678 3834
rect -644 3800 -608 3834
rect -574 3800 -538 3834
rect -504 3800 -468 3834
rect -434 3800 -398 3834
rect -364 3800 -328 3834
rect -271 3827 -258 3834
rect -197 3827 -188 3834
rect -123 3827 -118 3834
rect -294 3800 -258 3827
rect -224 3800 -188 3827
rect -154 3800 -118 3827
rect -84 3810 -48 3834
rect -14 3830 102 3834
rect -84 3800 -62 3810
rect -14 3800 68 3830
rect -852 3789 -62 3800
rect -852 3732 -818 3789
rect -784 3788 -62 3789
rect -784 3766 -305 3788
rect -271 3766 -231 3788
rect -197 3766 -157 3788
rect -123 3776 -62 3788
rect -28 3796 68 3800
rect -28 3776 102 3796
rect -123 3766 102 3776
rect -784 3732 -748 3766
rect -714 3732 -678 3766
rect -644 3732 -608 3766
rect -574 3732 -538 3766
rect -504 3732 -468 3766
rect -434 3732 -398 3766
rect -364 3732 -328 3766
rect -271 3754 -258 3766
rect -197 3754 -188 3766
rect -123 3754 -118 3766
rect -294 3732 -258 3754
rect -224 3732 -188 3754
rect -154 3732 -118 3754
rect -84 3738 -48 3766
rect -14 3762 102 3766
rect -84 3732 -62 3738
rect -14 3732 68 3762
rect -852 3717 -62 3732
rect -852 3664 -818 3717
rect -784 3715 -62 3717
rect -784 3698 -305 3715
rect -271 3698 -231 3715
rect -197 3698 -157 3715
rect -123 3704 -62 3715
rect -28 3728 68 3732
rect -28 3704 102 3728
rect -123 3698 102 3704
rect -784 3664 -748 3698
rect -714 3664 -678 3698
rect -644 3664 -608 3698
rect -574 3664 -538 3698
rect -504 3664 -468 3698
rect -434 3664 -398 3698
rect -364 3664 -328 3698
rect -271 3681 -258 3698
rect -197 3681 -188 3698
rect -123 3681 -118 3698
rect -294 3664 -258 3681
rect -224 3664 -188 3681
rect -154 3664 -118 3681
rect -84 3666 -48 3698
rect -14 3694 102 3698
rect -84 3664 -62 3666
rect -14 3664 68 3694
rect -852 3645 -62 3664
rect -852 3596 -818 3645
rect -784 3642 -62 3645
rect -784 3630 -305 3642
rect -271 3630 -231 3642
rect -197 3630 -157 3642
rect -123 3632 -62 3642
rect -28 3660 68 3664
rect -28 3632 102 3660
rect -123 3630 102 3632
rect -784 3596 -748 3630
rect -714 3596 -678 3630
rect -644 3596 -608 3630
rect -574 3596 -538 3630
rect -504 3596 -468 3630
rect -434 3596 -398 3630
rect -364 3596 -328 3630
rect -271 3608 -258 3630
rect -197 3608 -188 3630
rect -123 3608 -118 3630
rect -294 3596 -258 3608
rect -224 3596 -188 3608
rect -154 3596 -118 3608
rect -84 3596 -48 3630
rect -14 3626 102 3630
rect -14 3596 68 3626
rect -852 3594 68 3596
rect -852 3573 -62 3594
rect -852 3528 -818 3573
rect -784 3569 -62 3573
rect -784 3562 -305 3569
rect -271 3562 -231 3569
rect -197 3562 -157 3569
rect -123 3562 -62 3569
rect -28 3592 68 3594
rect -28 3562 102 3592
rect -784 3528 -748 3562
rect -714 3528 -678 3562
rect -644 3528 -608 3562
rect -574 3528 -538 3562
rect -504 3528 -468 3562
rect -434 3528 -398 3562
rect -364 3528 -328 3562
rect -271 3535 -258 3562
rect -197 3535 -188 3562
rect -123 3535 -118 3562
rect -294 3528 -258 3535
rect -224 3528 -188 3535
rect -154 3528 -118 3535
rect -84 3560 -62 3562
rect -84 3528 -48 3560
rect -14 3558 102 3562
rect -14 3528 68 3558
rect -852 3524 68 3528
rect -852 3522 102 3524
rect -852 3501 -62 3522
rect -852 3460 -818 3501
rect -784 3496 -62 3501
rect -784 3494 -305 3496
rect -271 3494 -231 3496
rect -197 3494 -157 3496
rect -123 3494 -62 3496
rect -28 3494 102 3522
rect -784 3460 -748 3494
rect -714 3460 -678 3494
rect -644 3460 -608 3494
rect -574 3460 -538 3494
rect -504 3460 -468 3494
rect -434 3460 -398 3494
rect -364 3460 -328 3494
rect -271 3462 -258 3494
rect -197 3462 -188 3494
rect -123 3462 -118 3494
rect -294 3460 -258 3462
rect -224 3460 -188 3462
rect -154 3460 -118 3462
rect -84 3488 -62 3494
rect -14 3490 102 3494
rect -84 3460 -48 3488
rect -14 3460 68 3490
rect -852 3456 68 3460
rect -852 3450 102 3456
rect -852 3429 -62 3450
rect -852 3392 -818 3429
rect -784 3426 -62 3429
rect -28 3426 102 3450
rect -784 3392 -748 3426
rect -714 3392 -678 3426
rect -644 3392 -608 3426
rect -574 3392 -538 3426
rect -504 3392 -468 3426
rect -434 3392 -398 3426
rect -364 3392 -328 3426
rect -294 3392 -258 3426
rect -224 3392 -188 3426
rect -154 3392 -118 3426
rect -84 3416 -62 3426
rect -14 3422 102 3426
rect -84 3392 -48 3416
rect -14 3392 68 3422
rect -852 3388 68 3392
rect -852 3378 102 3388
rect -852 3358 -62 3378
rect -28 3358 102 3378
rect -852 3323 -818 3358
rect -784 3324 -748 3358
rect -714 3324 -678 3358
rect -644 3324 -608 3358
rect -574 3324 -538 3358
rect -504 3324 -468 3358
rect -434 3324 -398 3358
rect -364 3324 -328 3358
rect -294 3324 -258 3358
rect -224 3324 -188 3358
rect -154 3324 -118 3358
rect -84 3344 -62 3358
rect -14 3354 102 3358
rect -84 3324 -48 3344
rect -14 3324 68 3354
rect -784 3323 68 3324
rect -852 3320 68 3323
rect -852 3306 102 3320
rect -852 3290 -62 3306
rect -28 3290 102 3306
rect -852 3251 -818 3290
rect -784 3256 -748 3290
rect -714 3256 -678 3290
rect -644 3256 -608 3290
rect -574 3256 -538 3290
rect -504 3256 -468 3290
rect -434 3256 -398 3290
rect -364 3256 -328 3290
rect -294 3256 -258 3290
rect -224 3256 -188 3290
rect -154 3256 -118 3290
rect -84 3272 -62 3290
rect -14 3286 102 3290
rect -84 3256 -48 3272
rect -14 3256 68 3286
rect -784 3252 68 3256
rect -784 3251 102 3252
rect -852 3234 102 3251
rect -852 3222 -62 3234
rect -28 3222 102 3234
rect -852 3179 -818 3222
rect -784 3188 -748 3222
rect -714 3188 -678 3222
rect -644 3188 -608 3222
rect -574 3188 -538 3222
rect -504 3188 -468 3222
rect -434 3188 -398 3222
rect -364 3188 -328 3222
rect -294 3188 -258 3222
rect -224 3188 -188 3222
rect -154 3188 -118 3222
rect -84 3200 -62 3222
rect -14 3218 102 3222
rect -84 3188 -48 3200
rect -14 3188 68 3218
rect -784 3184 68 3188
rect -784 3179 102 3184
rect -852 3154 102 3179
rect -852 3107 -818 3154
rect -784 3120 -748 3154
rect -714 3120 -678 3154
rect -644 3120 -608 3154
rect -574 3120 -538 3154
rect -504 3120 -468 3154
rect -434 3120 -398 3154
rect -364 3120 -328 3154
rect -294 3120 -258 3154
rect -224 3120 -188 3154
rect -154 3120 -118 3154
rect -84 3120 -48 3154
rect -14 3151 102 3154
rect -10 3150 102 3151
rect -784 3117 -44 3120
rect -10 3117 68 3150
rect -784 3116 68 3117
rect -784 3107 102 3116
rect -852 3086 102 3107
rect -852 3035 -818 3086
rect -784 3052 -748 3086
rect -714 3052 -678 3086
rect -644 3052 -608 3086
rect -574 3052 -538 3086
rect -504 3052 -468 3086
rect -434 3052 -398 3086
rect -364 3052 -328 3086
rect -294 3052 -258 3086
rect -224 3052 -188 3086
rect -154 3052 -118 3086
rect -84 3052 -48 3086
rect -14 3082 102 3086
rect -14 3079 68 3082
rect -784 3045 -44 3052
rect -10 3048 68 3079
rect -10 3045 102 3048
rect -784 3035 102 3045
rect -852 3018 102 3035
rect -852 2963 -818 3018
rect -784 2984 -748 3018
rect -714 2984 -678 3018
rect -644 2984 -608 3018
rect -574 2984 -538 3018
rect -504 2984 -468 3018
rect -434 2984 -398 3018
rect -364 2984 -328 3018
rect -294 2984 -258 3018
rect -224 2984 -188 3018
rect -154 2984 -118 3018
rect -84 2984 -48 3018
rect -14 3014 102 3018
rect -14 3007 68 3014
rect -784 2973 -44 2984
rect -10 2980 68 3007
rect -10 2973 102 2980
rect -784 2963 102 2973
rect -852 2950 102 2963
rect -852 2891 -818 2950
rect -784 2916 -748 2950
rect -714 2916 -678 2950
rect -644 2916 -608 2950
rect -574 2916 -538 2950
rect -504 2916 -468 2950
rect -434 2916 -398 2950
rect -364 2916 -328 2950
rect -294 2916 -258 2950
rect -224 2916 -188 2950
rect -154 2916 -118 2950
rect -84 2916 -48 2950
rect -14 2946 102 2950
rect -14 2935 68 2946
rect -784 2901 -44 2916
rect -10 2912 68 2935
rect -10 2901 102 2912
rect -784 2891 102 2901
rect -852 2882 102 2891
rect -852 2819 -818 2882
rect -784 2848 -748 2882
rect -714 2848 -678 2882
rect -644 2848 -608 2882
rect -574 2848 -538 2882
rect -504 2848 -468 2882
rect -434 2848 -398 2882
rect -364 2848 -328 2882
rect -294 2848 -258 2882
rect -224 2848 -188 2882
rect -154 2848 -118 2882
rect -84 2848 -48 2882
rect -14 2878 102 2882
rect -14 2863 68 2878
rect -784 2829 -44 2848
rect -10 2844 68 2863
rect -10 2829 102 2844
rect -784 2819 102 2829
rect -852 2814 102 2819
rect -852 2747 -818 2814
rect -784 2780 -748 2814
rect -714 2780 -678 2814
rect -644 2780 -608 2814
rect -574 2780 -538 2814
rect -504 2780 -468 2814
rect -434 2780 -398 2814
rect -364 2780 -328 2814
rect -294 2780 -258 2814
rect -224 2780 -188 2814
rect -154 2780 -118 2814
rect -84 2780 -48 2814
rect -14 2810 102 2814
rect -14 2791 68 2810
rect -784 2757 -44 2780
rect -10 2776 68 2791
rect -10 2757 102 2776
rect -784 2747 102 2757
rect -852 2746 102 2747
rect -852 2712 -818 2746
rect -784 2712 -748 2746
rect -714 2712 -678 2746
rect -644 2712 -608 2746
rect -574 2712 -538 2746
rect -504 2712 -468 2746
rect -434 2712 -398 2746
rect -364 2712 -328 2746
rect -294 2712 -258 2746
rect -224 2712 -188 2746
rect -154 2712 -118 2746
rect -84 2712 -48 2746
rect -14 2742 102 2746
rect -14 2719 68 2742
rect -852 2709 -44 2712
rect -852 2644 -818 2709
rect -784 2685 -44 2709
rect -10 2708 68 2719
rect -10 2685 102 2708
rect -784 2678 102 2685
rect -784 2644 -748 2678
rect -714 2644 -678 2678
rect -644 2644 -608 2678
rect -574 2644 -538 2678
rect -504 2644 -468 2678
rect -434 2644 -398 2678
rect -364 2644 -328 2678
rect -294 2644 -258 2678
rect -224 2644 -188 2678
rect -154 2644 -118 2678
rect -84 2644 -48 2678
rect -14 2674 102 2678
rect -14 2647 68 2674
rect -852 2637 -44 2644
rect -852 2576 -818 2637
rect -784 2613 -44 2637
rect -10 2640 68 2647
rect -10 2613 102 2640
rect -784 2610 102 2613
rect -784 2576 -748 2610
rect -714 2576 -678 2610
rect -644 2576 -608 2610
rect -574 2576 -538 2610
rect -504 2576 -468 2610
rect -434 2576 -398 2610
rect -364 2576 -328 2610
rect -294 2576 -258 2610
rect -224 2576 -188 2610
rect -154 2576 -118 2610
rect -84 2576 -48 2610
rect -14 2606 102 2610
rect -14 2576 68 2606
rect -852 2575 68 2576
rect -852 2565 -44 2575
rect -852 2508 -818 2565
rect -784 2542 -44 2565
rect -10 2572 68 2575
rect -784 2508 -748 2542
rect -714 2508 -678 2542
rect -644 2508 -608 2542
rect -574 2508 -538 2542
rect -504 2508 -468 2542
rect -434 2508 -398 2542
rect -364 2508 -328 2542
rect -294 2508 -258 2542
rect -224 2508 -188 2542
rect -154 2508 -118 2542
rect -84 2508 -48 2542
rect -10 2541 102 2572
rect -14 2538 102 2541
rect -14 2508 68 2538
rect -852 2504 68 2508
rect -852 2503 102 2504
rect -852 2493 -44 2503
rect -852 2439 -818 2493
rect -784 2473 -44 2493
rect -784 2439 -748 2473
rect -714 2439 -678 2473
rect -644 2439 -608 2473
rect -574 2439 -538 2473
rect -504 2439 -468 2473
rect -434 2439 -398 2473
rect -364 2439 -328 2473
rect -294 2439 -258 2473
rect -224 2439 -188 2473
rect -154 2439 -118 2473
rect -84 2439 -48 2473
rect -10 2470 102 2503
rect -10 2469 68 2470
rect -14 2439 68 2469
rect -852 2436 68 2439
rect -852 2431 102 2436
rect -852 2421 -44 2431
rect -852 2370 -818 2421
rect -784 2404 -44 2421
rect -784 2370 -748 2404
rect -714 2370 -678 2404
rect -644 2370 -608 2404
rect -574 2370 -538 2404
rect -504 2370 -468 2404
rect -434 2370 -398 2404
rect -364 2370 -328 2404
rect -294 2370 -258 2404
rect -224 2370 -188 2404
rect -154 2370 -118 2404
rect -84 2370 -48 2404
rect -10 2402 102 2431
rect -10 2397 68 2402
rect -14 2370 68 2397
rect -852 2368 68 2370
rect -852 2359 102 2368
rect -852 2349 -44 2359
rect -852 2301 -818 2349
rect -784 2335 -44 2349
rect -784 2301 -748 2335
rect -714 2301 -678 2335
rect -644 2301 -608 2335
rect -574 2301 -538 2335
rect -504 2301 -468 2335
rect -434 2301 -398 2335
rect -364 2301 -328 2335
rect -294 2301 -258 2335
rect -224 2301 -188 2335
rect -154 2301 -118 2335
rect -84 2301 -48 2335
rect -10 2334 102 2359
rect -10 2325 68 2334
rect -14 2301 68 2325
rect -852 2300 68 2301
rect -852 2287 102 2300
rect -852 2277 -44 2287
rect -852 2232 -818 2277
rect -784 2266 -44 2277
rect -10 2266 102 2287
rect -784 2232 -748 2266
rect -714 2232 -678 2266
rect -644 2232 -608 2266
rect -574 2232 -538 2266
rect -504 2232 -468 2266
rect -434 2232 -398 2266
rect -364 2232 -328 2266
rect -294 2232 -258 2266
rect -224 2232 -188 2266
rect -154 2232 -118 2266
rect -84 2232 -48 2266
rect -10 2253 68 2266
rect -14 2232 68 2253
rect -852 2215 102 2232
rect -852 2205 -44 2215
rect -852 2163 -818 2205
rect -784 2197 -44 2205
rect -10 2198 102 2215
rect -784 2163 -748 2197
rect -714 2163 -678 2197
rect -644 2163 -608 2197
rect -574 2163 -538 2197
rect -504 2163 -468 2197
rect -434 2163 -398 2197
rect -364 2163 -328 2197
rect -294 2163 -258 2197
rect -224 2163 -188 2197
rect -154 2163 -118 2197
rect -84 2163 -48 2197
rect -10 2181 68 2198
rect -14 2164 68 2181
rect -14 2163 102 2164
rect -852 2143 102 2163
rect -852 2133 -44 2143
rect -852 2094 -818 2133
rect -784 2128 -44 2133
rect -10 2130 102 2143
rect -784 2094 -748 2128
rect -714 2094 -678 2128
rect -644 2094 -608 2128
rect -574 2094 -538 2128
rect -504 2094 -468 2128
rect -434 2094 -398 2128
rect -364 2094 -328 2128
rect -294 2094 -258 2128
rect -224 2094 -188 2128
rect -154 2094 -118 2128
rect -84 2094 -48 2128
rect -10 2109 68 2130
rect -14 2096 68 2109
rect -14 2094 102 2096
rect -852 2071 102 2094
rect -852 2061 -44 2071
rect -852 2025 -818 2061
rect -784 2059 -44 2061
rect -10 2062 102 2071
rect -784 2025 -748 2059
rect -714 2025 -678 2059
rect -644 2025 -608 2059
rect -574 2025 -538 2059
rect -504 2025 -468 2059
rect -434 2025 -398 2059
rect -364 2025 -328 2059
rect -294 2025 -258 2059
rect -224 2025 -188 2059
rect -154 2025 -118 2059
rect -84 2025 -48 2059
rect -10 2037 68 2062
rect -14 2028 68 2037
rect -14 2025 102 2028
rect -852 1999 102 2025
rect -852 1990 -44 1999
rect -10 1994 102 1999
rect -852 1955 -818 1990
rect -784 1956 -748 1990
rect -714 1956 -678 1990
rect -644 1956 -608 1990
rect -574 1956 -538 1990
rect -504 1956 -468 1990
rect -434 1956 -398 1990
rect -364 1956 -328 1990
rect -294 1956 -258 1990
rect -224 1956 -188 1990
rect -154 1956 -118 1990
rect -84 1956 -48 1990
rect -10 1965 68 1994
rect -14 1960 68 1965
rect -14 1956 102 1960
rect -784 1955 102 1956
rect -852 1927 102 1955
rect -852 1921 -44 1927
rect -10 1926 102 1927
rect -852 1883 -818 1921
rect -784 1887 -748 1921
rect -714 1887 -678 1921
rect -644 1887 -608 1921
rect -574 1887 -538 1921
rect -504 1887 -468 1921
rect -434 1887 -398 1921
rect -364 1887 -328 1921
rect -294 1887 -258 1921
rect -224 1887 -188 1921
rect -154 1887 -118 1921
rect -84 1887 -48 1921
rect -10 1893 68 1926
rect -14 1892 68 1893
rect -14 1887 102 1892
rect -784 1883 102 1887
rect -852 1858 102 1883
rect -852 1855 68 1858
rect -852 1852 -44 1855
rect -852 1811 -818 1852
rect -784 1818 -748 1852
rect -714 1818 -678 1852
rect -644 1818 -608 1852
rect -574 1818 -538 1852
rect -504 1818 -468 1852
rect -434 1818 -398 1852
rect -364 1818 -328 1852
rect -294 1818 -258 1852
rect -224 1818 -188 1852
rect -154 1818 -118 1852
rect -84 1818 -48 1852
rect -10 1824 68 1855
rect -10 1821 102 1824
rect -14 1818 102 1821
rect -784 1811 102 1818
rect -852 1790 102 1811
rect -852 1783 68 1790
rect -852 1739 -818 1783
rect -784 1749 -748 1783
rect -714 1749 -678 1783
rect -644 1749 -608 1783
rect -574 1749 -538 1783
rect -504 1749 -468 1783
rect -434 1749 -398 1783
rect -364 1749 -328 1783
rect -294 1749 -258 1783
rect -224 1749 -188 1783
rect -154 1749 -118 1783
rect -84 1749 -48 1783
rect -10 1756 68 1783
rect -10 1749 102 1756
rect -784 1739 102 1749
rect -852 1722 102 1739
rect -852 1714 68 1722
rect -852 1667 -818 1714
rect -784 1680 -748 1714
rect -714 1680 -678 1714
rect -644 1680 -608 1714
rect -574 1680 -538 1714
rect -504 1680 -468 1714
rect -434 1680 -398 1714
rect -364 1680 -328 1714
rect -294 1680 -258 1714
rect -224 1680 -188 1714
rect -154 1680 -118 1714
rect -84 1680 -48 1714
rect -14 1711 68 1714
rect -10 1688 68 1711
rect -784 1677 -44 1680
rect -10 1677 102 1688
rect -784 1667 102 1677
rect -852 1654 102 1667
rect -852 1645 68 1654
rect -852 1595 -818 1645
rect -784 1611 -748 1645
rect -714 1611 -678 1645
rect -644 1611 -608 1645
rect -574 1611 -538 1645
rect -504 1611 -468 1645
rect -434 1611 -398 1645
rect -364 1611 -328 1645
rect -294 1611 -258 1645
rect -224 1611 -188 1645
rect -154 1611 -118 1645
rect -84 1611 -48 1645
rect -14 1639 68 1645
rect -10 1620 68 1639
rect -784 1605 -44 1611
rect -10 1605 102 1620
rect -784 1595 102 1605
rect -852 1586 102 1595
rect -852 1576 68 1586
rect -852 1523 -818 1576
rect -784 1542 -748 1576
rect -714 1542 -678 1576
rect -644 1542 -608 1576
rect -574 1542 -538 1576
rect -504 1542 -468 1576
rect -434 1542 -398 1576
rect -364 1542 -328 1576
rect -294 1542 -258 1576
rect -224 1542 -188 1576
rect -154 1542 -118 1576
rect -84 1542 -48 1576
rect -14 1567 68 1576
rect -10 1552 68 1567
rect -784 1533 -44 1542
rect -10 1533 102 1552
rect -784 1523 102 1533
rect -852 1518 102 1523
rect -852 1507 68 1518
rect -852 1451 -818 1507
rect -784 1473 -748 1507
rect -714 1473 -678 1507
rect -644 1473 -608 1507
rect -574 1473 -538 1507
rect -504 1473 -468 1507
rect -434 1473 -398 1507
rect -364 1473 -328 1507
rect -294 1473 -258 1507
rect -224 1473 -188 1507
rect -154 1473 -118 1507
rect -84 1473 -48 1507
rect -14 1495 68 1507
rect -10 1484 68 1495
rect -784 1461 -44 1473
rect -10 1461 102 1484
rect -784 1451 102 1461
rect -852 1450 102 1451
rect -852 1438 68 1450
rect -852 1379 -818 1438
rect -784 1404 -748 1438
rect -714 1404 -678 1438
rect -644 1404 -608 1438
rect -574 1404 -538 1438
rect -504 1404 -468 1438
rect -434 1404 -398 1438
rect -364 1404 -328 1438
rect -294 1404 -258 1438
rect -224 1404 -188 1438
rect -154 1404 -118 1438
rect -84 1404 -48 1438
rect -14 1423 68 1438
rect -10 1416 68 1423
rect -784 1389 -44 1404
rect -10 1389 102 1416
rect -784 1381 102 1389
rect -784 1379 68 1381
rect -852 1369 68 1379
rect -852 1307 -818 1369
rect -784 1335 -748 1369
rect -714 1335 -678 1369
rect -644 1335 -608 1369
rect -574 1335 -538 1369
rect -504 1335 -468 1369
rect -434 1335 -398 1369
rect -364 1335 -328 1369
rect -294 1335 -258 1369
rect -224 1335 -188 1369
rect -154 1335 -118 1369
rect -84 1335 -48 1369
rect -14 1351 68 1369
rect -10 1347 68 1351
rect -784 1317 -44 1335
rect -10 1317 102 1347
rect -784 1312 102 1317
rect -784 1307 68 1312
rect -852 1300 68 1307
rect -852 1235 -818 1300
rect -784 1266 -748 1300
rect -714 1266 -678 1300
rect -644 1266 -608 1300
rect -574 1266 -538 1300
rect -504 1266 -468 1300
rect -434 1266 -398 1300
rect -364 1266 -328 1300
rect -294 1266 -258 1300
rect -224 1266 -188 1300
rect -154 1266 -118 1300
rect -84 1266 -48 1300
rect -14 1279 68 1300
rect -10 1278 68 1279
rect -784 1245 -44 1266
rect -10 1245 102 1278
rect -784 1243 102 1245
rect -784 1235 68 1243
rect -852 1231 68 1235
rect -852 1163 -818 1231
rect -784 1197 -748 1231
rect -714 1197 -678 1231
rect -644 1197 -608 1231
rect -574 1197 -538 1231
rect -504 1197 -468 1231
rect -434 1197 -398 1231
rect -364 1197 -328 1231
rect -294 1197 -258 1231
rect -224 1197 -188 1231
rect -154 1197 -118 1231
rect -84 1197 -48 1231
rect -14 1209 68 1231
rect -14 1207 102 1209
rect -784 1173 -44 1197
rect -10 1174 102 1207
rect -10 1173 68 1174
rect -784 1163 68 1173
rect -852 1162 68 1163
rect -852 1128 -818 1162
rect -784 1128 -748 1162
rect -714 1128 -678 1162
rect -644 1128 -608 1162
rect -574 1128 -538 1162
rect -504 1128 -468 1162
rect -434 1128 -398 1162
rect -364 1128 -328 1162
rect -294 1128 -258 1162
rect -224 1128 -188 1162
rect -154 1128 -118 1162
rect -84 1128 -48 1162
rect -14 1140 68 1162
rect -14 1135 102 1140
rect -852 1125 -44 1128
rect -852 1059 -818 1125
rect -784 1101 -44 1125
rect -10 1105 102 1135
rect -10 1101 68 1105
rect -784 1093 68 1101
rect -784 1059 -748 1093
rect -714 1059 -678 1093
rect -644 1059 -608 1093
rect -574 1059 -538 1093
rect -504 1059 -468 1093
rect -434 1059 -398 1093
rect -364 1059 -328 1093
rect -294 1059 -258 1093
rect -224 1059 -188 1093
rect -154 1059 -118 1093
rect -84 1059 -48 1093
rect -14 1071 68 1093
rect -14 1063 102 1071
rect -852 1053 -44 1059
rect -852 990 -818 1053
rect -784 1029 -44 1053
rect -10 1036 102 1063
rect -10 1029 68 1036
rect -784 1024 68 1029
rect -784 990 -748 1024
rect -714 990 -678 1024
rect -644 990 -608 1024
rect -574 990 -538 1024
rect -504 990 -468 1024
rect -434 990 -398 1024
rect -364 990 -328 1024
rect -294 990 -258 1024
rect -224 990 -188 1024
rect -154 990 -118 1024
rect -84 990 -48 1024
rect -14 1002 68 1024
rect -14 990 102 1002
rect -852 981 -44 990
rect -852 921 -818 981
rect -784 956 -44 981
rect -10 967 102 990
rect -10 956 68 967
rect -784 955 68 956
rect -784 921 -748 955
rect -714 921 -678 955
rect -644 921 -608 955
rect -574 921 -538 955
rect -504 921 -468 955
rect -434 921 -398 955
rect -364 921 -328 955
rect -294 921 -258 955
rect -224 921 -188 955
rect -154 921 -118 955
rect -84 921 -48 955
rect -14 933 68 955
rect -14 921 102 933
rect -852 917 102 921
rect -852 909 -44 917
rect -852 852 -818 909
rect -784 886 -44 909
rect -10 898 102 917
rect -784 852 -748 886
rect -714 852 -678 886
rect -644 852 -608 886
rect -574 852 -538 886
rect -504 852 -468 886
rect -434 852 -398 886
rect -364 852 -328 886
rect -294 852 -258 886
rect -224 852 -188 886
rect -154 852 -118 886
rect -84 852 -48 886
rect -10 883 68 898
rect -14 864 68 883
rect -14 852 102 864
rect -852 844 102 852
rect -852 837 -44 844
rect -852 783 -818 837
rect -784 817 -44 837
rect -10 829 102 844
rect -784 783 -748 817
rect -714 783 -678 817
rect -644 783 -608 817
rect -574 783 -538 817
rect -504 783 -468 817
rect -434 783 -398 817
rect -364 783 -328 817
rect -294 783 -258 817
rect -224 783 -188 817
rect -154 783 -118 817
rect -84 783 -48 817
rect -10 810 68 829
rect -14 795 68 810
rect -14 783 102 795
rect -852 771 102 783
rect -852 765 -44 771
rect -852 714 -818 765
rect -784 748 -44 765
rect -10 760 102 771
rect -784 714 -748 748
rect -714 714 -678 748
rect -644 714 -608 748
rect -574 714 -538 748
rect -504 714 -468 748
rect -434 714 -398 748
rect -364 714 -328 748
rect -294 714 -258 748
rect -224 714 -188 748
rect -154 714 -118 748
rect -84 714 -48 748
rect -10 737 68 760
rect -14 726 68 737
rect -14 714 102 726
rect -852 698 102 714
rect -852 693 -44 698
rect -852 645 -818 693
rect -784 679 -44 693
rect -10 691 102 698
rect -784 645 -748 679
rect -714 645 -678 679
rect -644 645 -608 679
rect -574 645 -538 679
rect -504 645 -468 679
rect -434 645 -398 679
rect -364 645 -328 679
rect -294 645 -258 679
rect -224 645 -188 679
rect -154 645 -118 679
rect -84 645 -48 679
rect -10 664 68 691
rect -14 657 68 664
rect -14 645 102 657
rect -852 625 102 645
rect -852 621 -44 625
rect -852 576 -818 621
rect -784 610 -44 621
rect -10 622 102 625
rect -784 576 -748 610
rect -714 576 -678 610
rect -644 576 -608 610
rect -574 576 -538 610
rect -504 576 -468 610
rect -434 576 -398 610
rect -364 576 -328 610
rect -294 576 -258 610
rect -224 576 -188 610
rect -154 576 -118 610
rect -84 576 -48 610
rect -10 591 68 622
rect -14 588 68 591
rect -14 576 102 588
rect -852 553 102 576
rect -852 552 68 553
rect -852 548 -44 552
rect -852 507 -818 548
rect -784 541 -44 548
rect -784 507 -748 541
rect -714 507 -678 541
rect -644 507 -608 541
rect -574 507 -538 541
rect -504 507 -468 541
rect -434 507 -398 541
rect -364 507 -328 541
rect -294 507 -258 541
rect -224 507 -188 541
rect -154 507 -118 541
rect -84 507 -48 541
rect -10 519 68 552
rect -10 518 102 519
rect -14 507 102 518
rect -852 484 102 507
rect -852 479 68 484
rect -852 475 -44 479
rect -852 438 -818 475
rect -784 472 -44 475
rect -784 438 -748 472
rect -714 438 -678 472
rect -644 438 -608 472
rect -574 438 -538 472
rect -504 438 -468 472
rect -434 438 -398 472
rect -364 438 -328 472
rect -294 438 -258 472
rect -224 438 -188 472
rect -154 438 -118 472
rect -84 438 -48 472
rect -10 450 68 479
rect -10 445 102 450
rect -14 438 102 445
rect -852 415 102 438
rect -852 406 68 415
rect -852 403 -44 406
rect -852 368 -818 403
rect -784 369 -748 403
rect -714 369 -678 403
rect -644 369 -608 403
rect -574 369 -538 403
rect -504 369 -468 403
rect -434 369 -398 403
rect -364 369 -328 403
rect -294 369 -258 403
rect -224 369 -188 403
rect -154 369 -118 403
rect -84 369 -48 403
rect -10 381 68 406
rect -10 372 102 381
rect -14 369 102 372
rect -784 368 102 369
rect -852 346 102 368
rect -852 334 68 346
rect -852 295 -818 334
rect -784 300 -748 334
rect -714 300 -678 334
rect -644 300 -608 334
rect -574 300 -538 334
rect -504 300 -468 334
rect -434 300 -398 334
rect -364 300 -328 334
rect -294 300 -258 334
rect -224 300 -188 334
rect -154 300 -118 334
rect -84 300 -48 334
rect -14 333 68 334
rect -10 312 68 333
rect -784 299 -44 300
rect -10 299 102 312
rect -784 295 102 299
rect -852 277 102 295
rect -852 265 68 277
rect -852 222 -818 265
rect -784 231 -748 265
rect -714 231 -678 265
rect -644 231 -608 265
rect -574 231 -538 265
rect -504 231 -468 265
rect -434 231 -398 265
rect -364 231 -328 265
rect -294 231 -258 265
rect -224 231 -188 265
rect -154 231 -118 265
rect -84 231 -48 265
rect -14 260 68 265
rect -10 243 68 260
rect -784 226 -44 231
rect -10 226 102 243
rect -784 222 102 226
rect -852 208 102 222
rect -852 196 68 208
rect -852 149 -818 196
rect -784 162 -748 196
rect -714 162 -678 196
rect -644 162 -608 196
rect -574 162 -538 196
rect -504 162 -468 196
rect -434 162 -398 196
rect -364 162 -328 196
rect -294 162 -258 196
rect -224 162 -188 196
rect -154 162 -118 196
rect -84 162 -48 196
rect -14 187 68 196
rect -10 174 68 187
rect -784 153 -44 162
rect -10 153 102 174
rect 154 4842 796 4924
rect 154 4808 231 4842
rect 265 4822 303 4842
rect 265 4808 278 4822
rect 337 4808 375 4842
rect 409 4822 447 4842
rect 425 4808 447 4822
rect 481 4808 519 4842
rect 553 4822 796 4842
rect 154 4788 278 4808
rect 312 4788 391 4808
rect 425 4788 525 4808
rect 559 4798 796 4822
rect 559 4788 662 4798
rect 154 4782 662 4788
rect 154 4778 651 4782
rect 154 4744 171 4778
rect 205 4758 651 4778
rect 696 4764 796 4798
rect 205 4744 318 4758
rect 154 4728 318 4744
rect 154 4702 254 4728
rect 154 4668 171 4702
rect 205 4694 254 4702
rect 288 4694 318 4728
rect 523 4748 651 4758
rect 685 4748 796 4764
rect 523 4729 796 4748
rect 205 4668 318 4694
rect 154 4659 318 4668
rect 154 4626 254 4659
rect 288 4658 318 4659
rect 154 4592 171 4626
rect 205 4625 254 4626
rect 205 4624 284 4625
rect 205 4592 318 4624
rect 154 4590 318 4592
rect 154 4556 254 4590
rect 288 4583 318 4590
rect 154 4550 284 4556
rect 154 4516 171 4550
rect 205 4549 284 4550
rect 205 4521 318 4549
rect 205 4516 254 4521
rect 154 4487 254 4516
rect 288 4508 318 4521
rect 154 4474 284 4487
rect 154 4440 171 4474
rect 205 4452 318 4474
rect 205 4440 254 4452
rect 154 4418 254 4440
rect 288 4433 318 4452
rect 154 4399 284 4418
rect 154 4398 318 4399
rect 154 4364 171 4398
rect 205 4383 318 4398
rect 205 4364 254 4383
rect 154 4349 254 4364
rect 288 4357 318 4383
rect 154 4323 284 4349
rect 154 4322 318 4323
rect 154 4288 171 4322
rect 205 4314 318 4322
rect 205 4288 254 4314
rect 154 4280 254 4288
rect 288 4281 318 4314
rect 154 4247 284 4280
rect 154 4246 318 4247
rect 154 4212 171 4246
rect 205 4245 318 4246
rect 205 4212 254 4245
rect 154 4211 254 4212
rect 288 4211 318 4245
rect 154 4205 318 4211
rect 154 4176 284 4205
rect 154 4170 254 4176
rect 154 4136 171 4170
rect 205 4142 254 4170
rect 288 4142 318 4171
rect 205 4136 318 4142
rect 154 4129 318 4136
rect 154 4107 284 4129
rect 154 4093 254 4107
rect 154 4059 171 4093
rect 205 4073 254 4093
rect 288 4073 318 4095
rect 205 4059 318 4073
rect 154 4053 318 4059
rect 154 4038 284 4053
rect 154 4016 254 4038
rect 154 3982 171 4016
rect 205 4004 254 4016
rect 288 4004 318 4019
rect 205 3982 318 4004
rect 154 3977 318 3982
rect 154 3969 284 3977
rect 154 3939 254 3969
rect 154 3905 171 3939
rect 205 3935 254 3939
rect 288 3935 318 3943
rect 205 3905 318 3935
rect 154 3901 318 3905
rect 154 3900 284 3901
rect 154 3866 254 3900
rect 288 3866 318 3867
rect 154 3862 318 3866
rect 154 3828 171 3862
rect 205 3831 318 3862
rect 205 3828 254 3831
rect 154 3797 254 3828
rect 288 3825 318 3831
rect 154 3791 284 3797
rect 154 3785 318 3791
rect 154 3751 171 3785
rect 205 3762 318 3785
rect 205 3751 254 3762
rect 154 3728 254 3751
rect 288 3728 318 3762
rect 154 3708 318 3728
rect 154 3674 171 3708
rect 205 3693 318 3708
rect 205 3674 254 3693
rect 154 3659 254 3674
rect 288 3659 318 3693
rect 154 3631 318 3659
rect 154 3597 171 3631
rect 205 3624 318 3631
rect 205 3597 254 3624
rect 154 3590 254 3597
rect 288 3590 318 3624
rect 154 3555 318 3590
rect 154 3549 254 3555
rect 288 3549 318 3555
rect 154 3515 167 3549
rect 201 3521 254 3549
rect 201 3515 255 3521
rect 289 3515 318 3549
rect 154 3486 318 3515
rect 154 3476 254 3486
rect 154 3442 167 3476
rect 201 3452 254 3476
rect 288 3475 318 3486
rect 201 3442 255 3452
rect 154 3441 255 3442
rect 289 3441 318 3475
rect 154 3417 318 3441
rect 154 3404 254 3417
rect 154 3370 167 3404
rect 201 3383 254 3404
rect 288 3401 318 3417
rect 201 3370 255 3383
rect 154 3367 255 3370
rect 289 3367 318 3401
rect 154 3348 318 3367
rect 154 3332 254 3348
rect 154 3298 167 3332
rect 201 3314 254 3332
rect 288 3327 318 3348
rect 201 3298 255 3314
rect 154 3293 255 3298
rect 289 3293 318 3327
rect 154 3279 318 3293
rect 154 3260 254 3279
rect 154 3226 167 3260
rect 201 3245 254 3260
rect 288 3253 318 3279
rect 201 3226 255 3245
rect 154 3219 255 3226
rect 289 3219 318 3253
rect 154 3210 318 3219
rect 154 3188 254 3210
rect 154 3154 167 3188
rect 201 3176 254 3188
rect 288 3179 318 3210
rect 201 3154 255 3176
rect 154 3145 255 3154
rect 289 3145 318 3179
rect 154 3141 318 3145
rect 154 3116 254 3141
rect 154 3082 167 3116
rect 201 3107 254 3116
rect 288 3107 318 3141
rect 201 3105 318 3107
rect 201 3082 255 3105
rect 154 3072 255 3082
rect 154 3044 254 3072
rect 289 3071 318 3105
rect 154 3010 167 3044
rect 201 3038 254 3044
rect 288 3038 318 3071
rect 201 3031 318 3038
rect 201 3010 255 3031
rect 154 3003 255 3010
rect 154 2972 254 3003
rect 289 2997 318 3031
rect 154 2938 167 2972
rect 201 2969 254 2972
rect 288 2969 318 2997
rect 201 2957 318 2969
rect 201 2938 255 2957
rect 154 2934 255 2938
rect 154 2900 254 2934
rect 289 2923 318 2957
rect 288 2900 318 2923
rect 154 2866 167 2900
rect 201 2883 318 2900
rect 201 2866 255 2883
rect 154 2865 255 2866
rect 154 2831 254 2865
rect 289 2849 318 2883
rect 288 2831 318 2849
rect 154 2828 318 2831
rect 154 2794 167 2828
rect 201 2809 318 2828
rect 201 2796 255 2809
rect 201 2794 254 2796
rect 154 2762 254 2794
rect 289 2775 318 2809
rect 288 2762 318 2775
rect 154 2756 318 2762
rect 154 2722 167 2756
rect 201 2735 318 2756
rect 201 2727 255 2735
rect 201 2722 254 2727
rect 154 2693 254 2722
rect 289 2701 318 2735
rect 288 2693 318 2701
rect 154 2684 318 2693
rect 154 2650 167 2684
rect 201 2661 318 2684
rect 201 2658 255 2661
rect 201 2650 254 2658
rect 154 2624 254 2650
rect 289 2627 318 2661
rect 288 2624 318 2627
rect 154 2612 318 2624
rect 154 2578 167 2612
rect 201 2589 318 2612
rect 201 2578 254 2589
rect 288 2587 318 2589
rect 154 2555 254 2578
rect 154 2553 255 2555
rect 289 2553 318 2587
rect 154 2540 318 2553
rect 154 2506 167 2540
rect 201 2520 318 2540
rect 201 2506 254 2520
rect 288 2514 318 2520
rect 154 2486 254 2506
rect 154 2480 255 2486
rect 289 2480 318 2514
rect 154 2468 318 2480
rect 154 2434 167 2468
rect 201 2451 318 2468
rect 201 2434 254 2451
rect 288 2441 318 2451
rect 154 2417 254 2434
rect 154 2407 255 2417
rect 289 2407 318 2441
rect 154 2396 318 2407
rect 154 2362 167 2396
rect 201 2382 318 2396
rect 201 2362 254 2382
rect 288 2368 318 2382
rect 154 2348 254 2362
rect 154 2334 255 2348
rect 289 2334 318 2368
rect 154 2324 318 2334
rect 154 2290 167 2324
rect 201 2313 318 2324
rect 201 2290 254 2313
rect 288 2295 318 2313
rect 154 2279 254 2290
rect 154 2261 255 2279
rect 289 2261 318 2295
rect 154 2252 318 2261
rect 154 2218 167 2252
rect 201 2244 318 2252
rect 201 2218 254 2244
rect 288 2222 318 2244
rect 154 2210 254 2218
rect 154 2188 255 2210
rect 289 2188 318 2222
rect 154 2180 318 2188
rect 154 2146 167 2180
rect 201 2175 318 2180
rect 201 2146 254 2175
rect 288 2149 318 2175
rect 154 2141 254 2146
rect 154 2115 255 2141
rect 289 2115 318 2149
rect 154 2108 318 2115
rect 154 2074 167 2108
rect 201 2106 318 2108
rect 201 2074 254 2106
rect 288 2076 318 2106
rect 154 2072 254 2074
rect 154 2042 255 2072
rect 289 2042 318 2076
rect 154 2037 318 2042
rect 154 2036 254 2037
rect 154 2002 167 2036
rect 201 2003 254 2036
rect 288 2003 318 2037
rect 201 2002 255 2003
rect 154 1969 255 2002
rect 289 1969 318 2003
rect 154 1968 318 1969
rect 154 1964 254 1968
rect 154 1930 167 1964
rect 201 1934 254 1964
rect 288 1934 318 1968
rect 201 1930 318 1934
rect 154 1899 255 1930
rect 154 1892 254 1899
rect 289 1896 318 1930
rect 154 1858 167 1892
rect 201 1865 254 1892
rect 288 1865 318 1896
rect 201 1858 318 1865
rect 154 1857 318 1858
rect 154 1830 255 1857
rect 154 1820 254 1830
rect 289 1823 318 1857
rect 154 1786 167 1820
rect 201 1796 254 1820
rect 288 1796 318 1823
rect 201 1786 318 1796
rect 154 1784 318 1786
rect 154 1761 255 1784
rect 154 1748 254 1761
rect 289 1750 318 1784
rect 154 1714 167 1748
rect 201 1727 254 1748
rect 288 1727 318 1750
rect 201 1714 318 1727
rect 154 1711 318 1714
rect 154 1692 255 1711
rect 154 1676 254 1692
rect 289 1677 318 1711
rect 154 1642 167 1676
rect 201 1658 254 1676
rect 288 1658 318 1677
rect 201 1642 318 1658
rect 154 1638 318 1642
rect 154 1623 255 1638
rect 154 1604 254 1623
rect 289 1604 318 1638
rect 154 1570 167 1604
rect 201 1589 254 1604
rect 288 1589 318 1604
rect 201 1570 318 1589
rect 154 1565 318 1570
rect 154 1554 255 1565
rect 154 1532 254 1554
rect 154 1498 167 1532
rect 201 1520 254 1532
rect 289 1531 318 1565
rect 288 1520 318 1531
rect 201 1498 318 1520
rect 154 1492 318 1498
rect 154 1485 255 1492
rect 154 1460 254 1485
rect 154 1426 167 1460
rect 201 1451 254 1460
rect 289 1458 318 1492
rect 288 1451 318 1458
rect 201 1426 318 1451
rect 154 1419 318 1426
rect 154 1416 255 1419
rect 154 1388 254 1416
rect 154 1354 167 1388
rect 201 1382 254 1388
rect 289 1385 318 1419
rect 288 1382 318 1385
rect 201 1354 318 1382
rect 154 1347 318 1354
rect 154 1316 254 1347
rect 288 1346 318 1347
rect 154 1282 167 1316
rect 201 1313 254 1316
rect 201 1312 255 1313
rect 289 1312 318 1346
rect 201 1282 318 1312
rect 154 1278 318 1282
rect 154 1244 254 1278
rect 288 1273 318 1278
rect 154 1210 167 1244
rect 201 1239 255 1244
rect 289 1239 318 1273
rect 201 1210 318 1239
rect 154 1209 318 1210
rect 154 1175 254 1209
rect 288 1200 318 1209
rect 154 1172 255 1175
rect 154 1138 167 1172
rect 201 1166 255 1172
rect 289 1166 318 1200
rect 201 1140 318 1166
rect 201 1138 254 1140
rect 154 1106 254 1138
rect 288 1127 318 1140
rect 154 1100 255 1106
rect 154 1066 167 1100
rect 201 1093 255 1100
rect 289 1093 318 1127
rect 201 1071 318 1093
rect 201 1066 254 1071
rect 154 1037 254 1066
rect 288 1054 318 1071
rect 154 1028 255 1037
rect 154 994 167 1028
rect 201 1020 255 1028
rect 289 1020 318 1054
rect 201 1002 318 1020
rect 201 994 254 1002
rect 154 968 254 994
rect 288 981 318 1002
rect 154 956 255 968
rect 154 922 167 956
rect 201 947 255 956
rect 289 947 318 981
rect 201 933 318 947
rect 201 922 254 933
rect 154 899 254 922
rect 288 908 318 933
rect 154 884 255 899
rect 154 850 167 884
rect 201 874 255 884
rect 289 874 318 908
rect 201 864 318 874
rect 201 850 254 864
rect 154 830 254 850
rect 288 835 318 864
rect 154 812 255 830
rect 154 778 167 812
rect 201 801 255 812
rect 289 801 318 835
rect 201 795 318 801
rect 201 778 254 795
rect 154 761 254 778
rect 288 762 318 795
rect 154 740 255 761
rect 154 706 167 740
rect 201 728 255 740
rect 289 728 318 762
rect 201 726 318 728
rect 201 706 254 726
rect 154 692 254 706
rect 288 692 318 726
rect 154 689 318 692
rect 154 668 255 689
rect 154 634 167 668
rect 201 657 255 668
rect 201 634 254 657
rect 289 655 318 689
rect 154 623 254 634
rect 288 623 318 655
rect 154 616 318 623
rect 154 596 255 616
rect 154 562 167 596
rect 201 588 255 596
rect 201 562 254 588
rect 289 582 318 616
rect 154 554 254 562
rect 288 554 318 582
rect 154 543 318 554
rect 154 524 255 543
rect 154 490 167 524
rect 201 519 255 524
rect 201 490 254 519
rect 289 509 318 543
rect 154 485 254 490
rect 288 485 318 509
rect 154 470 318 485
rect 154 452 255 470
rect 154 418 167 452
rect 201 450 255 452
rect 201 418 254 450
rect 289 436 318 470
rect 154 416 254 418
rect 288 416 318 436
rect 154 397 318 416
rect 154 381 255 397
rect 154 380 254 381
rect 154 346 167 380
rect 201 347 254 380
rect 289 363 318 397
rect 288 347 318 363
rect 370 4702 471 4718
rect 404 4668 471 4702
rect 370 4634 471 4668
rect 404 4600 471 4634
rect 370 4566 471 4600
rect 404 4532 471 4566
rect 370 4498 471 4532
rect 404 4464 471 4498
rect 370 4430 471 4464
rect 404 4396 471 4430
rect 370 4362 471 4396
rect 404 4328 471 4362
rect 370 4294 471 4328
rect 404 4260 471 4294
rect 370 4226 471 4260
rect 404 4192 471 4226
rect 370 4158 471 4192
rect 404 4124 471 4158
rect 370 4090 471 4124
rect 404 4056 471 4090
rect 370 4022 471 4056
rect 404 3988 471 4022
rect 370 3954 471 3988
rect 404 3920 471 3954
rect 370 3886 471 3920
rect 404 3852 471 3886
rect 370 3818 471 3852
rect 404 3784 471 3818
rect 370 3725 471 3784
rect 523 4708 662 4729
rect 523 4702 651 4708
rect 523 4668 546 4702
rect 580 4674 651 4702
rect 696 4695 796 4729
rect 685 4674 796 4695
rect 580 4668 796 4674
rect 523 4660 796 4668
rect 523 4658 662 4660
rect 523 4624 539 4658
rect 573 4634 662 4658
rect 523 4600 546 4624
rect 580 4600 651 4634
rect 696 4626 796 4660
rect 685 4600 796 4626
rect 523 4591 796 4600
rect 523 4583 662 4591
rect 523 4549 539 4583
rect 573 4566 662 4583
rect 580 4561 662 4566
rect 523 4532 546 4549
rect 580 4532 651 4561
rect 696 4557 796 4591
rect 523 4527 651 4532
rect 685 4527 796 4557
rect 523 4522 796 4527
rect 523 4508 662 4522
rect 523 4474 539 4508
rect 573 4498 662 4508
rect 580 4488 662 4498
rect 696 4488 796 4522
rect 523 4464 546 4474
rect 580 4464 651 4488
rect 523 4454 651 4464
rect 685 4454 796 4488
rect 523 4453 796 4454
rect 523 4433 662 4453
rect 523 4399 539 4433
rect 573 4430 662 4433
rect 580 4419 662 4430
rect 696 4419 796 4453
rect 580 4415 796 4419
rect 523 4396 546 4399
rect 580 4396 651 4415
rect 523 4381 651 4396
rect 685 4384 796 4415
rect 523 4362 662 4381
rect 523 4357 546 4362
rect 523 4323 539 4357
rect 580 4350 662 4362
rect 696 4350 796 4384
rect 580 4342 796 4350
rect 580 4328 651 4342
rect 573 4323 651 4328
rect 523 4308 651 4323
rect 685 4315 796 4342
rect 523 4294 662 4308
rect 523 4281 546 4294
rect 580 4281 662 4294
rect 696 4281 796 4315
rect 523 4247 539 4281
rect 580 4269 796 4281
rect 580 4260 651 4269
rect 573 4247 651 4260
rect 523 4235 651 4247
rect 685 4246 796 4269
rect 523 4226 662 4235
rect 523 4205 546 4226
rect 580 4212 662 4226
rect 696 4212 796 4246
rect 523 4171 539 4205
rect 580 4196 796 4212
rect 580 4192 651 4196
rect 573 4171 651 4192
rect 685 4177 796 4196
rect 523 4162 651 4171
rect 523 4158 662 4162
rect 523 4129 546 4158
rect 580 4143 662 4158
rect 696 4143 796 4177
rect 523 4095 539 4129
rect 580 4124 796 4143
rect 573 4123 796 4124
rect 573 4095 651 4123
rect 685 4108 796 4123
rect 523 4090 651 4095
rect 523 4056 546 4090
rect 580 4089 651 4090
rect 580 4074 662 4089
rect 696 4074 796 4108
rect 580 4056 796 4074
rect 523 4053 796 4056
rect 523 4019 539 4053
rect 573 4050 796 4053
rect 573 4022 651 4050
rect 685 4039 796 4050
rect 523 3988 546 4019
rect 580 4016 651 4022
rect 580 4005 662 4016
rect 696 4005 796 4039
rect 580 3988 796 4005
rect 523 3977 796 3988
rect 523 3943 539 3977
rect 573 3954 651 3977
rect 685 3970 796 3977
rect 580 3943 651 3954
rect 523 3920 546 3943
rect 580 3936 662 3943
rect 696 3936 796 3970
rect 580 3920 796 3936
rect 523 3904 796 3920
rect 523 3901 651 3904
rect 685 3901 796 3904
rect 523 3867 539 3901
rect 573 3886 651 3901
rect 580 3870 651 3886
rect 580 3867 662 3870
rect 696 3867 796 3901
rect 523 3852 546 3867
rect 580 3852 796 3867
rect 523 3832 796 3852
rect 523 3831 662 3832
rect 523 3825 651 3831
rect 523 3791 539 3825
rect 573 3818 651 3825
rect 580 3797 651 3818
rect 696 3798 796 3832
rect 685 3797 796 3798
rect 523 3784 546 3791
rect 580 3784 796 3797
rect 523 3763 796 3784
rect 523 3758 662 3763
rect 523 3725 651 3758
rect 696 3729 796 3763
rect 370 3694 438 3725
rect 404 3660 438 3694
rect 546 3724 651 3725
rect 685 3724 796 3729
rect 546 3694 796 3724
rect 370 3621 438 3660
rect 404 3587 438 3621
rect 370 3581 438 3587
rect 404 3514 438 3581
rect 370 3513 438 3514
rect 404 3479 438 3513
rect 370 3475 438 3479
rect 404 3411 438 3475
rect 370 3402 438 3411
rect 404 3343 438 3402
rect 370 3329 438 3343
rect 404 3275 438 3329
rect 370 3256 438 3275
rect 404 3207 438 3256
rect 370 3183 438 3207
rect 404 3139 438 3183
rect 370 3110 438 3139
rect 404 3071 438 3110
rect 370 3037 438 3071
rect 404 3003 438 3037
rect 370 2969 438 3003
rect 404 2930 438 2969
rect 370 2901 438 2930
rect 404 2857 438 2901
rect 370 2833 438 2857
rect 404 2784 438 2833
rect 370 2765 438 2784
rect 404 2711 438 2765
rect 370 2697 438 2711
rect 404 2639 438 2697
rect 370 2601 438 2639
rect 404 2567 438 2601
rect 370 2529 438 2567
rect 404 2495 438 2529
rect 370 2460 438 2495
rect 404 2423 438 2460
rect 370 2392 438 2423
rect 404 2351 438 2392
rect 370 2324 438 2351
rect 404 2279 438 2324
rect 370 2256 438 2279
rect 404 2207 438 2256
rect 370 2188 438 2207
rect 404 2135 438 2188
rect 370 2120 438 2135
rect 404 2063 438 2120
rect 370 2052 438 2063
rect 404 2018 438 2052
rect 370 2016 438 2018
rect 404 1950 438 2016
rect 370 1943 438 1950
rect 404 1882 438 1943
rect 370 1870 438 1882
rect 404 1814 438 1870
rect 370 1797 438 1814
rect 404 1746 438 1797
rect 370 1725 438 1746
rect 404 1678 438 1725
rect 370 1653 438 1678
rect 404 1610 438 1653
rect 370 1581 438 1610
rect 404 1542 438 1581
rect 370 1509 438 1542
rect 404 1475 438 1509
rect 370 1437 438 1475
rect 404 1403 438 1437
rect 370 1365 438 1403
rect 472 3674 506 3690
rect 472 3586 506 3625
rect 472 3513 506 3552
rect 472 3440 506 3479
rect 472 3367 506 3406
rect 472 3294 506 3333
rect 472 3221 506 3260
rect 472 3148 506 3187
rect 472 3074 506 3114
rect 472 3000 506 3040
rect 472 2926 506 2966
rect 472 2852 506 2892
rect 472 2778 506 2818
rect 472 2704 506 2744
rect 472 2630 506 2670
rect 472 2556 506 2596
rect 472 2482 506 2519
rect 472 2408 506 2448
rect 472 2334 506 2374
rect 472 2260 506 2300
rect 472 2186 506 2226
rect 472 2112 506 2152
rect 472 2038 506 2078
rect 472 1964 506 2004
rect 472 1890 506 1930
rect 472 1816 506 1856
rect 472 1742 506 1782
rect 472 1668 506 1708
rect 472 1594 506 1634
rect 472 1520 506 1560
rect 472 1446 506 1486
rect 472 1384 506 1400
rect 546 3685 662 3694
rect 546 3651 651 3685
rect 696 3660 796 3694
rect 685 3651 796 3660
rect 546 3625 796 3651
rect 546 3612 662 3625
rect 546 3581 651 3612
rect 696 3591 796 3625
rect 580 3578 651 3581
rect 685 3578 796 3591
rect 580 3556 796 3578
rect 580 3547 662 3556
rect 546 3539 662 3547
rect 546 3513 651 3539
rect 696 3522 796 3556
rect 580 3505 651 3513
rect 685 3505 796 3522
rect 580 3487 796 3505
rect 580 3479 662 3487
rect 546 3466 662 3479
rect 546 3445 651 3466
rect 696 3453 796 3487
rect 580 3432 651 3445
rect 685 3432 796 3453
rect 580 3418 796 3432
rect 580 3411 662 3418
rect 546 3393 662 3411
rect 546 3377 651 3393
rect 696 3384 796 3418
rect 580 3359 651 3377
rect 685 3359 796 3384
rect 580 3349 796 3359
rect 580 3343 662 3349
rect 546 3320 662 3343
rect 546 3309 651 3320
rect 696 3315 796 3349
rect 580 3286 651 3309
rect 685 3286 796 3315
rect 580 3280 796 3286
rect 580 3275 662 3280
rect 546 3247 662 3275
rect 546 3241 651 3247
rect 696 3246 796 3280
rect 580 3213 651 3241
rect 685 3213 796 3246
rect 580 3211 796 3213
rect 580 3207 662 3211
rect 546 3177 662 3207
rect 696 3177 796 3211
rect 546 3174 796 3177
rect 546 3173 651 3174
rect 580 3140 651 3173
rect 685 3142 796 3174
rect 580 3139 662 3140
rect 546 3108 662 3139
rect 696 3108 796 3142
rect 546 3105 796 3108
rect 580 3101 796 3105
rect 580 3071 651 3101
rect 685 3073 796 3101
rect 546 3067 651 3071
rect 546 3039 662 3067
rect 696 3039 796 3073
rect 546 3037 796 3039
rect 580 3028 796 3037
rect 580 3003 651 3028
rect 685 3004 796 3028
rect 546 2994 651 3003
rect 546 2970 662 2994
rect 696 2970 796 3004
rect 546 2969 796 2970
rect 580 2955 796 2969
rect 580 2935 651 2955
rect 685 2935 796 2955
rect 546 2921 651 2935
rect 546 2901 662 2921
rect 696 2901 796 2935
rect 580 2882 796 2901
rect 580 2867 651 2882
rect 546 2848 651 2867
rect 685 2866 796 2882
rect 546 2833 662 2848
rect 580 2832 662 2833
rect 696 2832 796 2866
rect 580 2809 796 2832
rect 580 2799 651 2809
rect 546 2775 651 2799
rect 685 2797 796 2809
rect 546 2765 662 2775
rect 580 2763 662 2765
rect 696 2763 796 2797
rect 580 2736 796 2763
rect 580 2731 651 2736
rect 546 2702 651 2731
rect 685 2728 796 2736
rect 546 2697 662 2702
rect 580 2694 662 2697
rect 696 2694 796 2728
rect 580 2663 796 2694
rect 546 2629 651 2663
rect 685 2659 796 2663
rect 546 2625 662 2629
rect 696 2625 796 2659
rect 546 2590 796 2625
rect 546 2556 651 2590
rect 696 2556 796 2590
rect 546 2521 796 2556
rect 546 2517 662 2521
rect 546 2483 651 2517
rect 696 2487 796 2521
rect 685 2483 796 2487
rect 546 2460 796 2483
rect 580 2452 796 2460
rect 580 2444 662 2452
rect 580 2426 651 2444
rect 546 2410 651 2426
rect 696 2418 796 2452
rect 685 2410 796 2418
rect 546 2392 796 2410
rect 580 2383 796 2392
rect 580 2371 662 2383
rect 580 2358 651 2371
rect 546 2337 651 2358
rect 696 2349 796 2383
rect 685 2337 796 2349
rect 546 2324 796 2337
rect 580 2314 796 2324
rect 580 2298 662 2314
rect 580 2290 651 2298
rect 546 2264 651 2290
rect 696 2280 796 2314
rect 685 2264 796 2280
rect 546 2256 796 2264
rect 580 2245 796 2256
rect 580 2225 662 2245
rect 580 2222 651 2225
rect 546 2191 651 2222
rect 696 2211 796 2245
rect 685 2191 796 2211
rect 546 2188 796 2191
rect 580 2176 796 2188
rect 580 2154 662 2176
rect 546 2152 662 2154
rect 546 2120 651 2152
rect 696 2142 796 2176
rect 580 2118 651 2120
rect 685 2118 796 2142
rect 580 2107 796 2118
rect 580 2086 662 2107
rect 546 2079 662 2086
rect 546 2052 651 2079
rect 696 2073 796 2107
rect 580 2045 651 2052
rect 685 2045 796 2073
rect 580 2038 796 2045
rect 580 2018 662 2038
rect 546 2004 662 2018
rect 696 2004 796 2038
rect 546 1984 796 2004
rect 580 1969 796 1984
rect 580 1950 662 1969
rect 546 1935 662 1950
rect 696 1935 796 1969
rect 546 1924 796 1935
rect 546 1916 668 1924
rect 580 1900 668 1916
rect 580 1882 662 1900
rect 702 1890 756 1924
rect 790 1890 796 1924
rect 546 1866 662 1882
rect 696 1866 796 1890
rect 546 1852 796 1866
rect 546 1848 668 1852
rect 580 1831 668 1848
rect 702 1851 796 1852
rect 580 1814 662 1831
rect 702 1818 756 1851
rect 546 1797 662 1814
rect 696 1817 756 1818
rect 790 1817 796 1851
rect 696 1797 796 1817
rect 546 1780 796 1797
rect 580 1762 668 1780
rect 702 1778 796 1780
rect 580 1746 662 1762
rect 702 1746 756 1778
rect 546 1728 662 1746
rect 696 1744 756 1746
rect 790 1744 796 1778
rect 696 1728 796 1744
rect 546 1712 796 1728
rect 580 1708 796 1712
rect 580 1693 668 1708
rect 702 1705 796 1708
rect 580 1678 662 1693
rect 546 1659 662 1678
rect 702 1674 756 1705
rect 696 1671 756 1674
rect 790 1671 796 1705
rect 696 1659 796 1671
rect 546 1644 796 1659
rect 580 1636 796 1644
rect 580 1624 668 1636
rect 702 1632 796 1636
rect 580 1610 662 1624
rect 546 1590 662 1610
rect 702 1602 756 1632
rect 696 1598 756 1602
rect 790 1598 796 1632
rect 696 1590 796 1598
rect 546 1576 796 1590
rect 580 1564 796 1576
rect 580 1555 668 1564
rect 702 1559 796 1564
rect 580 1542 662 1555
rect 546 1521 662 1542
rect 702 1530 756 1559
rect 696 1525 756 1530
rect 790 1525 796 1559
rect 696 1521 796 1525
rect 546 1492 796 1521
rect 546 1486 668 1492
rect 702 1486 796 1492
rect 546 1452 662 1486
rect 702 1458 756 1486
rect 696 1452 756 1458
rect 790 1452 796 1486
rect 546 1419 796 1452
rect 546 1417 668 1419
rect 404 1344 438 1365
rect 546 1383 662 1417
rect 702 1413 796 1419
rect 702 1385 756 1413
rect 696 1383 756 1385
rect 546 1379 756 1383
rect 790 1379 796 1413
rect 546 1348 796 1379
rect 546 1344 662 1348
rect 696 1346 796 1348
rect 404 1331 471 1344
rect 370 1293 471 1331
rect 404 1258 471 1293
rect 370 1224 471 1258
rect 404 1187 471 1224
rect 370 1156 471 1187
rect 404 1115 471 1156
rect 370 1088 471 1115
rect 404 1043 471 1088
rect 370 1020 471 1043
rect 404 971 471 1020
rect 370 952 471 971
rect 404 899 471 952
rect 370 884 471 899
rect 404 827 471 884
rect 370 816 471 827
rect 404 755 471 816
rect 370 748 471 755
rect 404 683 471 748
rect 370 680 471 683
rect 404 646 471 680
rect 370 645 471 646
rect 404 578 471 645
rect 370 573 471 578
rect 404 510 471 573
rect 370 501 471 510
rect 404 442 471 501
rect 370 408 471 442
rect 404 374 471 408
rect 370 358 471 374
rect 523 1314 662 1344
rect 702 1340 796 1346
rect 523 1312 668 1314
rect 702 1312 756 1340
rect 523 1306 756 1312
rect 790 1306 796 1340
rect 523 1292 796 1306
rect 523 1258 546 1292
rect 580 1279 796 1292
rect 580 1258 662 1279
rect 696 1273 796 1279
rect 523 1245 662 1258
rect 702 1267 796 1273
rect 523 1239 668 1245
rect 702 1239 756 1267
rect 523 1233 756 1239
rect 790 1233 796 1267
rect 523 1224 796 1233
rect 523 1190 546 1224
rect 580 1210 796 1224
rect 580 1190 662 1210
rect 696 1200 796 1210
rect 523 1176 662 1190
rect 702 1194 796 1200
rect 523 1166 668 1176
rect 702 1166 756 1194
rect 523 1160 756 1166
rect 790 1160 796 1194
rect 523 1156 796 1160
rect 523 1122 546 1156
rect 580 1141 796 1156
rect 580 1122 662 1141
rect 696 1127 796 1141
rect 523 1107 662 1122
rect 702 1121 796 1127
rect 523 1093 668 1107
rect 702 1093 756 1121
rect 523 1088 756 1093
rect 523 1054 546 1088
rect 580 1087 756 1088
rect 790 1087 796 1121
rect 580 1072 796 1087
rect 580 1054 662 1072
rect 696 1054 796 1072
rect 523 1038 662 1054
rect 702 1048 796 1054
rect 523 1020 668 1038
rect 702 1020 756 1048
rect 523 986 546 1020
rect 580 1014 756 1020
rect 790 1014 796 1048
rect 580 1003 796 1014
rect 580 986 662 1003
rect 523 969 662 986
rect 696 981 796 1003
rect 702 974 796 981
rect 523 952 668 969
rect 523 918 546 952
rect 580 947 668 952
rect 702 947 756 974
rect 580 940 756 947
rect 790 940 796 974
rect 580 934 796 940
rect 580 918 662 934
rect 523 900 662 918
rect 696 908 796 934
rect 702 900 796 908
rect 523 884 668 900
rect 523 850 546 884
rect 580 874 668 884
rect 702 874 756 900
rect 580 866 756 874
rect 790 866 796 900
rect 580 865 796 866
rect 580 850 662 865
rect 523 831 662 850
rect 696 835 796 865
rect 523 816 668 831
rect 523 782 546 816
rect 580 801 668 816
rect 702 826 796 835
rect 702 801 756 826
rect 580 796 756 801
rect 580 782 662 796
rect 523 762 662 782
rect 696 792 756 796
rect 790 792 796 826
rect 696 762 796 792
rect 523 748 668 762
rect 523 714 546 748
rect 580 728 668 748
rect 702 752 796 762
rect 702 728 756 752
rect 580 727 756 728
rect 580 714 662 727
rect 523 693 662 714
rect 696 718 756 727
rect 790 718 796 752
rect 696 693 796 718
rect 523 689 796 693
rect 523 680 668 689
rect 523 646 546 680
rect 580 658 668 680
rect 702 678 796 689
rect 580 646 662 658
rect 702 655 756 678
rect 523 624 662 646
rect 696 644 756 655
rect 790 644 796 678
rect 696 624 796 644
rect 523 616 796 624
rect 523 612 668 616
rect 523 578 546 612
rect 580 589 668 612
rect 702 604 796 616
rect 580 578 662 589
rect 702 582 756 604
rect 523 555 662 578
rect 696 570 756 582
rect 790 570 796 604
rect 696 555 796 570
rect 523 544 796 555
rect 523 510 546 544
rect 580 543 796 544
rect 580 520 668 543
rect 702 530 796 543
rect 580 510 662 520
rect 523 486 662 510
rect 702 509 756 530
rect 696 496 756 509
rect 790 496 796 530
rect 696 486 796 496
rect 523 476 796 486
rect 523 442 546 476
rect 580 470 796 476
rect 580 451 668 470
rect 702 456 796 470
rect 580 442 662 451
rect 523 417 662 442
rect 702 436 756 456
rect 696 422 756 436
rect 790 422 796 456
rect 696 417 796 422
rect 523 408 796 417
rect 523 374 546 408
rect 580 397 796 408
rect 580 382 668 397
rect 702 382 796 397
rect 580 374 662 382
rect 201 346 318 347
rect 154 324 318 346
rect 523 348 662 374
rect 702 363 756 382
rect 696 348 756 363
rect 790 348 796 382
rect 523 324 796 348
rect 154 312 255 324
rect 154 308 254 312
rect 154 274 167 308
rect 201 278 254 308
rect 289 290 338 324
rect 372 290 421 324
rect 455 290 504 324
rect 538 290 586 324
rect 620 290 668 324
rect 702 308 796 324
rect 702 290 756 308
rect 288 288 756 290
rect 288 278 352 288
rect 201 274 352 278
rect 154 254 352 274
rect 386 254 423 288
rect 457 254 494 288
rect 528 254 566 288
rect 600 254 638 288
rect 672 274 756 288
rect 790 274 796 308
rect 672 254 796 274
rect 154 236 796 254
rect 154 202 239 236
rect 273 202 313 236
rect 347 202 387 236
rect 421 202 461 236
rect 495 202 535 236
rect 569 202 609 236
rect 643 202 683 236
rect 717 202 796 236
rect 154 154 796 202
rect -784 149 102 153
rect -852 127 102 149
rect -852 76 -818 127
rect -784 93 -748 127
rect -714 93 -678 127
rect -644 93 -608 127
rect -574 93 -538 127
rect -504 93 -468 127
rect -434 93 -398 127
rect -364 93 -328 127
rect -294 93 -258 127
rect -224 93 -188 127
rect -154 93 -118 127
rect -84 93 -48 127
rect -14 114 102 127
rect -10 102 102 114
rect 848 102 882 4976
rect -10 95 92 102
rect 126 95 161 102
rect 195 95 230 102
rect 264 95 300 102
rect 334 95 370 102
rect 404 95 440 102
rect 474 95 510 102
rect -784 80 -44 93
rect -10 80 59 95
rect -784 76 59 80
rect -852 61 59 76
rect 126 68 134 95
rect 195 68 209 95
rect 264 68 284 95
rect 334 68 359 95
rect 404 68 434 95
rect 474 68 509 95
rect 544 68 580 102
rect 614 95 650 102
rect 684 95 720 102
rect 754 95 790 102
rect 824 95 882 102
rect 618 68 650 95
rect 693 68 720 95
rect 768 68 790 95
rect 93 61 134 68
rect 168 61 209 68
rect 243 61 284 68
rect 318 61 359 68
rect 393 61 434 68
rect 468 61 509 68
rect 543 61 584 68
rect 618 61 659 68
rect 693 61 734 68
rect 768 61 808 68
rect 842 61 882 95
rect -852 58 882 61
rect -852 3 -818 58
rect -784 24 -748 58
rect -714 24 -678 58
rect -644 24 -608 58
rect -574 24 -538 58
rect -504 24 -468 58
rect -434 24 -398 58
rect -364 24 -328 58
rect -294 24 -258 58
rect -224 24 -188 58
rect -154 24 -118 58
rect -84 24 -48 58
rect -14 41 882 58
rect -10 34 882 41
rect -784 7 -44 24
rect -10 19 92 34
rect 126 19 161 34
rect 195 19 230 34
rect -10 7 36 19
rect -784 3 36 7
rect -852 -15 36 3
rect 70 0 92 19
rect 147 0 161 19
rect 224 0 230 19
rect 264 19 300 34
rect 334 19 370 34
rect 404 19 440 34
rect 474 19 510 34
rect 544 19 580 34
rect 264 0 267 19
rect 334 0 344 19
rect 404 0 421 19
rect 474 0 498 19
rect 544 0 575 19
rect 614 0 650 34
rect 684 19 720 34
rect 754 19 790 34
rect 824 19 882 34
rect 687 0 720 19
rect 765 0 790 19
rect 70 -15 113 0
rect 147 -15 190 0
rect 224 -15 267 0
rect 301 -15 344 0
rect 378 -15 421 0
rect 455 -15 498 0
rect 532 -15 575 0
rect 609 -15 653 0
rect 687 -15 731 0
rect 765 -15 809 0
rect 843 -15 882 19
rect -852 -33 882 -15
rect -852 -34 898 -33
rect -852 -70 -818 -34
rect -784 -68 -750 -34
rect -716 -68 -682 -34
rect -648 -68 -614 -34
rect -580 -68 -546 -34
rect -512 -68 -478 -34
rect -444 -68 -410 -34
rect -376 -68 -342 -34
rect -308 -68 -274 -34
rect -240 -68 -205 -34
rect -171 -68 -136 -34
rect -102 -68 -67 -34
rect -33 -68 2 -34
rect 36 -65 71 -34
rect -784 -70 36 -68
rect -852 -99 36 -70
rect 70 -68 71 -65
rect 105 -65 140 -34
rect 174 -65 209 -34
rect 243 -65 278 -34
rect 312 -65 347 -34
rect 105 -68 113 -65
rect 174 -68 190 -65
rect 243 -68 267 -65
rect 312 -68 344 -65
rect 381 -68 416 -34
rect 450 -65 485 -34
rect 519 -65 554 -34
rect 588 -65 623 -34
rect 657 -65 692 -34
rect 455 -68 485 -65
rect 532 -68 554 -65
rect 609 -68 623 -65
rect 687 -68 692 -65
rect 726 -65 761 -34
rect 795 -65 830 -34
rect 726 -68 731 -65
rect 795 -68 809 -65
rect 864 -68 898 -34
rect 70 -99 113 -68
rect 147 -99 190 -68
rect 224 -99 267 -68
rect 301 -99 344 -68
rect 378 -99 421 -68
rect 455 -99 498 -68
rect 532 -99 575 -68
rect 609 -99 653 -68
rect 687 -99 731 -68
rect 765 -99 809 -68
rect 843 -99 898 -68
rect -852 -105 898 -99
rect -852 -143 -818 -105
rect -784 -139 -750 -105
rect -716 -139 -682 -105
rect -648 -139 -614 -105
rect -580 -139 -546 -105
rect -512 -139 -478 -105
rect -444 -139 -410 -105
rect -376 -139 -342 -105
rect -308 -139 -274 -105
rect -240 -139 -205 -105
rect -171 -139 -136 -105
rect -102 -139 -67 -105
rect -33 -139 2 -105
rect 36 -139 71 -105
rect 105 -139 140 -105
rect 174 -139 209 -105
rect 243 -139 278 -105
rect 312 -139 347 -105
rect 381 -139 416 -105
rect 450 -139 485 -105
rect 519 -139 554 -105
rect 588 -139 623 -105
rect 657 -139 692 -105
rect 726 -139 761 -105
rect 795 -139 830 -105
rect 864 -139 898 -105
rect -784 -143 898 -139
rect -852 -149 898 -143
rect -852 -176 36 -149
rect -852 -216 -818 -176
rect -784 -210 -750 -176
rect -716 -210 -682 -176
rect -648 -210 -614 -176
rect -580 -210 -546 -176
rect -512 -210 -478 -176
rect -444 -210 -410 -176
rect -376 -210 -342 -176
rect -308 -210 -274 -176
rect -240 -210 -205 -176
rect -171 -210 -136 -176
rect -102 -210 -67 -176
rect -33 -210 2 -176
rect 70 -176 113 -149
rect 147 -176 190 -149
rect 224 -176 267 -149
rect 301 -176 344 -149
rect 378 -176 421 -149
rect 455 -176 498 -149
rect 532 -176 575 -149
rect 609 -176 653 -149
rect 687 -176 731 -149
rect 765 -176 809 -149
rect 843 -176 898 -149
rect 70 -183 71 -176
rect 36 -210 71 -183
rect 105 -183 113 -176
rect 174 -183 190 -176
rect 243 -183 267 -176
rect 312 -183 344 -176
rect 105 -210 140 -183
rect 174 -210 209 -183
rect 243 -210 278 -183
rect 312 -210 347 -183
rect 381 -210 416 -176
rect 455 -183 485 -176
rect 532 -183 554 -176
rect 609 -183 623 -176
rect 687 -183 692 -176
rect 450 -210 485 -183
rect 519 -210 554 -183
rect 588 -210 623 -183
rect 657 -210 692 -183
rect 726 -183 731 -176
rect 795 -183 809 -176
rect 726 -210 761 -183
rect 795 -210 830 -183
rect 864 -210 898 -176
rect -784 -215 898 -210
rect -784 -216 -42 -215
rect -852 -247 -42 -216
rect -8 -233 898 -215
rect -8 -247 36 -233
rect -852 -289 -818 -247
rect -784 -281 -750 -247
rect -716 -255 -682 -247
rect -696 -281 -682 -255
rect -648 -281 -614 -247
rect -580 -281 -546 -247
rect -512 -281 -478 -247
rect -444 -281 -410 -247
rect -376 -281 -342 -247
rect -308 -281 -274 -247
rect -240 -281 -205 -247
rect -171 -281 -136 -247
rect -102 -281 -67 -247
rect -8 -249 2 -247
rect -33 -281 2 -249
rect 70 -247 113 -233
rect 147 -247 190 -233
rect 224 -247 267 -233
rect 301 -247 344 -233
rect 378 -247 421 -233
rect 455 -247 498 -233
rect 532 -247 575 -233
rect 609 -247 653 -233
rect 687 -247 731 -233
rect 765 -247 809 -233
rect 843 -247 898 -233
rect 70 -267 71 -247
rect 36 -281 71 -267
rect 105 -267 113 -247
rect 174 -267 190 -247
rect 243 -267 267 -247
rect 312 -267 344 -247
rect 105 -281 140 -267
rect 174 -281 209 -267
rect 243 -281 278 -267
rect 312 -281 347 -267
rect 381 -281 416 -247
rect 455 -267 485 -247
rect 532 -267 554 -247
rect 609 -267 623 -247
rect 687 -267 692 -247
rect 450 -281 485 -267
rect 519 -281 554 -267
rect 588 -281 623 -267
rect 657 -281 692 -267
rect 726 -267 731 -247
rect 795 -267 809 -247
rect 726 -281 761 -267
rect 795 -281 830 -267
rect 864 -281 898 -247
rect -784 -289 -730 -281
rect -696 -287 898 -281
rect -696 -289 -114 -287
rect -852 -318 -114 -289
rect -80 -318 -42 -287
rect -8 -317 898 -287
rect -8 -318 36 -317
rect -852 -352 -818 -318
rect -784 -352 -750 -318
rect -716 -327 -682 -318
rect -696 -352 -682 -327
rect -648 -352 -614 -318
rect -580 -352 -546 -318
rect -512 -352 -478 -318
rect -444 -352 -410 -318
rect -376 -352 -342 -318
rect -308 -352 -274 -318
rect -240 -352 -205 -318
rect -171 -352 -136 -318
rect -80 -321 -67 -318
rect -8 -321 2 -318
rect -102 -352 -67 -321
rect -33 -352 2 -321
rect 70 -318 113 -317
rect 147 -318 190 -317
rect 224 -318 267 -317
rect 301 -318 344 -317
rect 378 -318 421 -317
rect 455 -318 498 -317
rect 532 -318 575 -317
rect 609 -318 653 -317
rect 687 -318 731 -317
rect 765 -318 809 -317
rect 843 -318 898 -317
rect 70 -351 71 -318
rect 36 -352 71 -351
rect 105 -351 113 -318
rect 174 -351 190 -318
rect 243 -351 267 -318
rect 312 -351 344 -318
rect 105 -352 140 -351
rect 174 -352 209 -351
rect 243 -352 278 -351
rect 312 -352 347 -351
rect 381 -352 416 -318
rect 455 -351 485 -318
rect 532 -351 554 -318
rect 609 -351 623 -318
rect 687 -351 692 -318
rect 450 -352 485 -351
rect 519 -352 554 -351
rect 588 -352 623 -351
rect 657 -352 692 -351
rect 726 -351 731 -318
rect 795 -351 809 -318
rect 726 -352 761 -351
rect 795 -352 830 -351
rect 864 -352 898 -318
rect -852 -353 -730 -352
rect -696 -353 898 -352
rect 36 -354 843 -353
<< viali >>
rect -818 14504 -794 14517
rect -794 14504 -784 14517
rect -305 14504 -276 14505
rect -276 14504 -271 14505
rect -231 14504 -207 14505
rect -207 14504 -197 14505
rect -157 14504 -138 14505
rect -138 14504 -123 14505
rect -818 14483 -784 14504
rect -305 14471 -271 14504
rect -231 14471 -197 14504
rect -157 14471 -123 14504
rect -818 14432 -794 14445
rect -794 14432 -784 14445
rect -305 14432 -276 14433
rect -276 14432 -271 14433
rect -231 14432 -207 14433
rect -207 14432 -197 14433
rect -157 14432 -138 14433
rect -138 14432 -123 14433
rect 211 14432 241 14462
rect 241 14432 245 14462
rect 293 14432 310 14462
rect 310 14432 327 14462
rect 375 14432 379 14462
rect 379 14432 409 14462
rect 457 14432 483 14462
rect 483 14432 491 14462
rect 539 14432 552 14462
rect 552 14432 573 14462
rect 621 14432 655 14462
rect 703 14432 724 14462
rect 724 14432 737 14462
rect -818 14411 -784 14432
rect -305 14399 -271 14432
rect -231 14399 -197 14432
rect -157 14399 -123 14432
rect 211 14428 245 14432
rect 293 14428 327 14432
rect 375 14428 409 14432
rect 457 14428 491 14432
rect 539 14428 573 14432
rect 621 14428 655 14432
rect 703 14428 737 14432
rect -818 14360 -794 14373
rect -794 14360 -784 14373
rect -305 14360 -276 14361
rect -276 14360 -271 14361
rect -231 14360 -207 14361
rect -207 14360 -197 14361
rect -157 14360 -138 14361
rect -138 14360 -123 14361
rect 211 14360 241 14389
rect 241 14360 245 14389
rect 293 14360 310 14389
rect 310 14360 327 14389
rect 375 14360 379 14389
rect 379 14360 409 14389
rect 457 14360 483 14389
rect 483 14360 491 14389
rect 539 14360 552 14389
rect 552 14360 573 14389
rect 621 14360 655 14389
rect 703 14360 724 14389
rect 724 14360 737 14389
rect -818 14339 -784 14360
rect -305 14327 -271 14360
rect -231 14327 -197 14360
rect -157 14327 -123 14360
rect 211 14355 245 14360
rect 293 14355 327 14360
rect 375 14355 409 14360
rect 457 14355 491 14360
rect 539 14355 573 14360
rect 621 14355 655 14360
rect 703 14355 737 14360
rect -818 14288 -794 14301
rect -794 14288 -784 14301
rect -305 14288 -276 14289
rect -276 14288 -271 14289
rect -231 14288 -207 14289
rect -207 14288 -197 14289
rect -157 14288 -138 14289
rect -138 14288 -123 14289
rect 211 14288 241 14316
rect 241 14288 245 14316
rect 293 14288 310 14316
rect 310 14288 327 14316
rect 375 14288 379 14316
rect 379 14288 409 14316
rect 457 14288 483 14316
rect 483 14288 491 14316
rect 539 14288 552 14316
rect 552 14288 573 14316
rect 621 14288 655 14316
rect 703 14288 724 14316
rect 724 14288 737 14316
rect -818 14267 -784 14288
rect -305 14255 -271 14288
rect -231 14255 -197 14288
rect -157 14255 -123 14288
rect 211 14282 245 14288
rect 293 14282 327 14288
rect 375 14282 409 14288
rect 457 14282 491 14288
rect 539 14282 573 14288
rect 621 14282 655 14288
rect 703 14282 737 14288
rect -818 14216 -794 14229
rect -794 14216 -784 14229
rect -305 14216 -276 14217
rect -276 14216 -271 14217
rect -231 14216 -207 14217
rect -207 14216 -197 14217
rect -157 14216 -138 14217
rect -138 14216 -123 14217
rect 211 14216 241 14243
rect 241 14216 245 14243
rect 293 14216 310 14243
rect 310 14216 327 14243
rect 375 14216 379 14243
rect 379 14216 409 14243
rect 457 14216 483 14243
rect 483 14216 491 14243
rect 539 14216 552 14243
rect 552 14216 573 14243
rect 621 14216 655 14243
rect 703 14216 724 14243
rect 724 14216 737 14243
rect -818 14195 -784 14216
rect -305 14183 -271 14216
rect -231 14183 -197 14216
rect -157 14183 -123 14216
rect 211 14209 245 14216
rect 293 14209 327 14216
rect 375 14209 409 14216
rect 457 14209 491 14216
rect 539 14209 573 14216
rect 621 14209 655 14216
rect 703 14209 737 14216
rect -818 14144 -794 14157
rect -794 14144 -784 14157
rect -305 14144 -276 14145
rect -276 14144 -271 14145
rect -231 14144 -207 14145
rect -207 14144 -197 14145
rect -157 14144 -138 14145
rect -138 14144 -123 14145
rect 211 14144 241 14170
rect 241 14144 245 14170
rect 293 14144 310 14170
rect 310 14144 327 14170
rect 375 14144 379 14170
rect 379 14144 409 14170
rect 457 14144 483 14170
rect 483 14144 491 14170
rect 539 14144 552 14170
rect 552 14144 573 14170
rect 621 14144 655 14170
rect 703 14144 724 14170
rect 724 14144 737 14170
rect -818 14123 -784 14144
rect -305 14111 -271 14144
rect -231 14111 -197 14144
rect -157 14111 -123 14144
rect 211 14136 245 14144
rect 293 14136 327 14144
rect 375 14136 409 14144
rect 457 14136 491 14144
rect 539 14136 573 14144
rect 621 14136 655 14144
rect 703 14136 737 14144
rect -818 14072 -794 14085
rect -794 14072 -784 14085
rect -305 14072 -276 14073
rect -276 14072 -271 14073
rect -231 14072 -207 14073
rect -207 14072 -197 14073
rect -157 14072 -138 14073
rect -138 14072 -123 14073
rect 211 14072 241 14097
rect 241 14072 245 14097
rect 293 14072 310 14097
rect 310 14072 327 14097
rect 375 14072 379 14097
rect 379 14072 409 14097
rect 457 14072 483 14097
rect 483 14072 491 14097
rect 539 14072 552 14097
rect 552 14072 573 14097
rect 621 14072 655 14097
rect 703 14072 724 14097
rect 724 14072 737 14097
rect -818 14051 -784 14072
rect -305 14039 -271 14072
rect -231 14039 -197 14072
rect -157 14039 -123 14072
rect 211 14063 245 14072
rect 293 14063 327 14072
rect 375 14063 409 14072
rect 457 14063 491 14072
rect 539 14063 573 14072
rect 621 14063 655 14072
rect 703 14063 737 14072
rect -818 14000 -794 14013
rect -794 14000 -784 14013
rect -305 14000 -276 14001
rect -276 14000 -271 14001
rect -231 14000 -207 14001
rect -207 14000 -197 14001
rect -157 14000 -138 14001
rect -138 14000 -123 14001
rect 211 14000 241 14024
rect 241 14000 245 14024
rect 293 14000 310 14024
rect 310 14000 327 14024
rect 375 14000 379 14024
rect 379 14000 409 14024
rect 457 14000 483 14024
rect 483 14000 491 14024
rect 539 14000 552 14024
rect 552 14000 573 14024
rect 621 14000 655 14024
rect 703 14000 724 14024
rect 724 14000 737 14024
rect -818 13979 -784 14000
rect -305 13967 -271 14000
rect -231 13967 -197 14000
rect -157 13967 -123 14000
rect -818 13932 -784 13941
rect -818 13907 -784 13932
rect -305 13898 -271 13929
rect -231 13898 -197 13929
rect -157 13898 -123 13929
rect -818 13864 -784 13869
rect -305 13895 -294 13898
rect -294 13895 -271 13898
rect -231 13895 -224 13898
rect -224 13895 -197 13898
rect -157 13895 -154 13898
rect -154 13895 -123 13898
rect -818 13835 -784 13864
rect -305 13830 -271 13857
rect -231 13830 -197 13857
rect -157 13830 -123 13857
rect -818 13796 -784 13797
rect -305 13823 -294 13830
rect -294 13823 -271 13830
rect -231 13823 -224 13830
rect -224 13823 -197 13830
rect -157 13823 -154 13830
rect -154 13823 -123 13830
rect -818 13763 -784 13796
rect -305 13762 -271 13785
rect -231 13762 -197 13785
rect -157 13762 -123 13785
rect -305 13751 -294 13762
rect -294 13751 -271 13762
rect -231 13751 -224 13762
rect -224 13751 -197 13762
rect -157 13751 -154 13762
rect -154 13751 -123 13762
rect -818 13694 -784 13725
rect -305 13694 -271 13713
rect -231 13694 -197 13713
rect -157 13694 -123 13713
rect -818 13691 -784 13694
rect -305 13679 -294 13694
rect -294 13679 -271 13694
rect -231 13679 -224 13694
rect -224 13679 -197 13694
rect -157 13679 -154 13694
rect -154 13679 -123 13694
rect -818 13626 -784 13653
rect -305 13626 -271 13641
rect -231 13626 -197 13641
rect -157 13626 -123 13641
rect -818 13619 -784 13626
rect -305 13607 -294 13626
rect -294 13607 -271 13626
rect -231 13607 -224 13626
rect -224 13607 -197 13626
rect -157 13607 -154 13626
rect -154 13607 -123 13626
rect -818 13558 -784 13581
rect -305 13558 -271 13569
rect -231 13558 -197 13569
rect -157 13558 -123 13569
rect -818 13547 -784 13558
rect -305 13535 -294 13558
rect -294 13535 -271 13558
rect -231 13535 -224 13558
rect -224 13535 -197 13558
rect -157 13535 -154 13558
rect -154 13535 -123 13558
rect -818 13490 -784 13509
rect -305 13490 -271 13497
rect -231 13490 -197 13497
rect -157 13490 -123 13497
rect -818 13475 -784 13490
rect -305 13463 -294 13490
rect -294 13463 -271 13490
rect -231 13463 -224 13490
rect -224 13463 -197 13490
rect -157 13463 -154 13490
rect -154 13463 -123 13490
rect -818 13422 -784 13437
rect -305 13422 -271 13425
rect -231 13422 -197 13425
rect -157 13422 -123 13425
rect -818 13403 -784 13422
rect -305 13391 -294 13422
rect -294 13391 -271 13422
rect -231 13391 -224 13422
rect -224 13391 -197 13422
rect -157 13391 -154 13422
rect -154 13391 -123 13422
rect -818 13354 -784 13365
rect -818 13331 -784 13354
rect -305 13320 -294 13353
rect -294 13320 -271 13353
rect -231 13320 -224 13353
rect -224 13320 -197 13353
rect -157 13320 -154 13353
rect -154 13320 -123 13353
rect -305 13319 -271 13320
rect -231 13319 -197 13320
rect -157 13319 -123 13320
rect -818 13286 -784 13293
rect -818 13259 -784 13286
rect -305 13252 -294 13281
rect -294 13252 -271 13281
rect -231 13252 -224 13281
rect -224 13252 -197 13281
rect -157 13252 -154 13281
rect -154 13252 -123 13281
rect -305 13247 -271 13252
rect -231 13247 -197 13252
rect -157 13247 -123 13252
rect -818 13218 -784 13221
rect -818 13187 -784 13218
rect -305 13184 -294 13209
rect -294 13184 -271 13209
rect -231 13184 -224 13209
rect -224 13184 -197 13209
rect -157 13184 -154 13209
rect -154 13184 -123 13209
rect -305 13175 -271 13184
rect -231 13175 -197 13184
rect -157 13175 -123 13184
rect -818 13116 -784 13149
rect -305 13116 -294 13137
rect -294 13116 -271 13137
rect -231 13116 -224 13137
rect -224 13116 -197 13137
rect -157 13116 -154 13137
rect -154 13116 -123 13137
rect -818 13115 -784 13116
rect -305 13103 -271 13116
rect -231 13103 -197 13116
rect -157 13103 -123 13116
rect -818 13048 -784 13077
rect -305 13048 -294 13065
rect -294 13048 -271 13065
rect -231 13048 -224 13065
rect -224 13048 -197 13065
rect -157 13048 -154 13065
rect -154 13048 -123 13065
rect -818 13043 -784 13048
rect -305 13031 -271 13048
rect -231 13031 -197 13048
rect -157 13031 -123 13048
rect -818 12980 -784 13005
rect -305 12980 -294 12993
rect -294 12980 -271 12993
rect -231 12980 -224 12993
rect -224 12980 -197 12993
rect -157 12980 -154 12993
rect -154 12980 -123 12993
rect -818 12971 -784 12980
rect -305 12959 -271 12980
rect -231 12959 -197 12980
rect -157 12959 -123 12980
rect -818 12912 -784 12933
rect -305 12912 -294 12921
rect -294 12912 -271 12921
rect -231 12912 -224 12921
rect -224 12912 -197 12921
rect -157 12912 -154 12921
rect -154 12912 -123 12921
rect -818 12899 -784 12912
rect -305 12887 -271 12912
rect -231 12887 -197 12912
rect -157 12887 -123 12912
rect -818 12844 -784 12861
rect -305 12844 -294 12849
rect -294 12844 -271 12849
rect -231 12844 -224 12849
rect -224 12844 -197 12849
rect -157 12844 -154 12849
rect -154 12844 -123 12849
rect -818 12827 -784 12844
rect -305 12815 -271 12844
rect -231 12815 -197 12844
rect -157 12815 -123 12844
rect -818 12776 -784 12789
rect -305 12776 -294 12777
rect -294 12776 -271 12777
rect -231 12776 -224 12777
rect -224 12776 -197 12777
rect -157 12776 -154 12777
rect -154 12776 -123 12777
rect -818 12755 -784 12776
rect -305 12743 -271 12776
rect -231 12743 -197 12776
rect -157 12743 -123 12776
rect -818 12708 -784 12717
rect -818 12683 -784 12708
rect -305 12674 -271 12705
rect -231 12674 -197 12705
rect -157 12674 -123 12705
rect -818 12640 -784 12645
rect -305 12671 -294 12674
rect -294 12671 -271 12674
rect -231 12671 -224 12674
rect -224 12671 -197 12674
rect -157 12671 -154 12674
rect -154 12671 -123 12674
rect -818 12611 -784 12640
rect -305 12606 -271 12633
rect -231 12606 -197 12633
rect -157 12606 -123 12633
rect -818 12572 -784 12573
rect -305 12599 -294 12606
rect -294 12599 -271 12606
rect -231 12599 -224 12606
rect -224 12599 -197 12606
rect -157 12599 -154 12606
rect -154 12599 -123 12606
rect -818 12539 -784 12572
rect -305 12538 -271 12561
rect -231 12538 -197 12561
rect -157 12538 -123 12561
rect -305 12527 -294 12538
rect -294 12527 -271 12538
rect -231 12527 -224 12538
rect -224 12527 -197 12538
rect -157 12527 -154 12538
rect -154 12527 -123 12538
rect -818 12470 -784 12501
rect -305 12470 -271 12489
rect -231 12470 -197 12489
rect -157 12470 -123 12489
rect -818 12467 -784 12470
rect -305 12455 -294 12470
rect -294 12455 -271 12470
rect -231 12455 -224 12470
rect -224 12455 -197 12470
rect -157 12455 -154 12470
rect -154 12455 -123 12470
rect 211 13990 245 14000
rect 293 13990 327 14000
rect 375 13990 409 14000
rect 457 13990 491 14000
rect 539 13990 573 14000
rect 621 13990 655 14000
rect 703 13990 737 14000
rect 211 13917 245 13951
rect 293 13917 327 13951
rect 375 13917 409 13951
rect 457 13917 491 13951
rect 539 13917 573 13951
rect 621 13917 655 13951
rect 703 13917 737 13951
rect 211 13844 245 13878
rect 293 13844 327 13878
rect 375 13844 409 13878
rect 457 13844 491 13878
rect 539 13844 573 13878
rect 621 13844 655 13878
rect 703 13844 737 13878
rect 211 13771 245 13805
rect 293 13771 327 13805
rect 375 13771 409 13805
rect 457 13771 491 13805
rect 539 13771 573 13805
rect 621 13771 655 13805
rect 703 13771 737 13805
rect 211 13698 245 13732
rect 293 13698 327 13732
rect 375 13698 409 13732
rect 457 13698 491 13732
rect 539 13698 573 13732
rect 621 13698 655 13732
rect 703 13698 737 13732
rect 211 13624 245 13658
rect 293 13624 327 13658
rect 375 13624 409 13658
rect 457 13624 491 13658
rect 539 13624 573 13658
rect 621 13624 655 13658
rect 703 13624 737 13658
rect 211 13550 245 13584
rect 293 13550 327 13584
rect 375 13550 409 13584
rect 457 13550 491 13584
rect 539 13550 573 13584
rect 621 13550 655 13584
rect 703 13550 737 13584
rect 211 13476 245 13510
rect 293 13476 327 13510
rect 375 13476 409 13510
rect 457 13476 491 13510
rect 539 13476 573 13510
rect 621 13476 655 13510
rect 703 13476 737 13510
rect 211 13402 245 13436
rect 293 13402 327 13436
rect 375 13402 409 13436
rect 457 13402 491 13436
rect 539 13402 573 13436
rect 621 13402 655 13436
rect 703 13402 737 13436
rect 211 13328 245 13362
rect 293 13328 327 13362
rect 375 13328 409 13362
rect 457 13328 491 13362
rect 539 13328 573 13362
rect 621 13328 655 13362
rect 703 13328 737 13362
rect 211 13254 245 13288
rect 293 13254 327 13288
rect 375 13254 409 13288
rect 457 13254 491 13288
rect 539 13254 573 13288
rect 621 13254 655 13288
rect 703 13254 737 13288
rect 211 13180 245 13214
rect 293 13180 327 13214
rect 375 13180 409 13214
rect 457 13180 491 13214
rect 539 13180 573 13214
rect 621 13180 655 13214
rect 703 13180 737 13214
rect 211 13106 245 13140
rect 293 13106 327 13140
rect 375 13106 409 13140
rect 457 13106 491 13140
rect 539 13106 573 13140
rect 621 13106 655 13140
rect 703 13106 737 13140
rect 211 13032 245 13066
rect 293 13032 327 13066
rect 375 13032 409 13066
rect 457 13032 491 13066
rect 539 13032 573 13066
rect 621 13032 655 13066
rect 703 13032 737 13066
rect 211 12958 245 12992
rect 293 12958 327 12992
rect 375 12958 409 12992
rect 457 12958 491 12992
rect 539 12958 573 12992
rect 621 12958 655 12992
rect 703 12958 737 12992
rect 211 12884 245 12918
rect 293 12884 327 12918
rect 375 12884 409 12918
rect 457 12884 491 12918
rect 539 12884 573 12918
rect 621 12884 655 12918
rect 703 12884 737 12918
rect 211 12810 245 12844
rect 293 12810 327 12844
rect 375 12810 409 12844
rect 457 12810 491 12844
rect 539 12810 573 12844
rect 621 12810 655 12844
rect 703 12810 737 12844
rect 211 12736 245 12770
rect 293 12736 327 12770
rect 375 12736 409 12770
rect 457 12736 491 12770
rect 539 12736 573 12770
rect 621 12736 655 12770
rect 703 12736 737 12770
rect 211 12662 245 12696
rect 293 12662 327 12696
rect 375 12662 409 12696
rect 457 12662 491 12696
rect 539 12662 573 12696
rect 621 12662 655 12696
rect 703 12662 737 12696
rect 211 12588 245 12622
rect 293 12588 327 12622
rect 375 12588 409 12622
rect 457 12588 491 12622
rect 539 12588 573 12622
rect 621 12588 655 12622
rect 703 12588 737 12622
rect 211 12514 245 12548
rect 293 12514 327 12548
rect 375 12514 409 12548
rect 457 12514 491 12548
rect 539 12514 573 12548
rect 621 12514 655 12548
rect 703 12514 737 12548
rect 211 12440 245 12474
rect 293 12440 327 12474
rect 375 12440 409 12474
rect 457 12440 491 12474
rect 539 12440 573 12474
rect 621 12440 655 12474
rect 703 12440 737 12474
rect -818 12402 -784 12429
rect -305 12402 -271 12417
rect -231 12402 -197 12417
rect -157 12402 -123 12417
rect -818 12395 -784 12402
rect -305 12383 -294 12402
rect -294 12383 -271 12402
rect -231 12383 -224 12402
rect -224 12383 -197 12402
rect -157 12383 -154 12402
rect -154 12383 -123 12402
rect -818 12334 -784 12357
rect -305 12334 -271 12345
rect -231 12334 -197 12345
rect -157 12334 -123 12345
rect -818 12323 -784 12334
rect -305 12311 -294 12334
rect -294 12311 -271 12334
rect -231 12311 -224 12334
rect -224 12311 -197 12334
rect -157 12311 -154 12334
rect -154 12311 -123 12334
rect -818 12266 -784 12285
rect -305 12266 -271 12273
rect -231 12266 -197 12273
rect -157 12266 -123 12273
rect -818 12251 -784 12266
rect -305 12239 -294 12266
rect -294 12239 -271 12266
rect -231 12239 -224 12266
rect -224 12239 -197 12266
rect -157 12239 -154 12266
rect -154 12239 -123 12266
rect -818 12198 -784 12213
rect -305 12198 -271 12201
rect -231 12198 -197 12201
rect -157 12198 -123 12201
rect -818 12179 -784 12198
rect -305 12167 -294 12198
rect -294 12167 -271 12198
rect -231 12167 -224 12198
rect -224 12167 -197 12198
rect -157 12167 -154 12198
rect -154 12167 -123 12198
rect -818 12130 -784 12141
rect -818 12107 -784 12130
rect -305 12096 -294 12129
rect -294 12096 -271 12129
rect -231 12096 -224 12129
rect -224 12096 -197 12129
rect -157 12096 -154 12129
rect -154 12096 -123 12129
rect -305 12095 -271 12096
rect -231 12095 -197 12096
rect -157 12095 -123 12096
rect -818 12062 -784 12069
rect -818 12035 -784 12062
rect -305 12028 -294 12057
rect -294 12028 -271 12057
rect -231 12028 -224 12057
rect -224 12028 -197 12057
rect -157 12028 -154 12057
rect -154 12028 -123 12057
rect -305 12023 -271 12028
rect -231 12023 -197 12028
rect -157 12023 -123 12028
rect -818 11994 -784 11997
rect -818 11963 -784 11994
rect -305 11960 -294 11985
rect -294 11960 -271 11985
rect -231 11960 -224 11985
rect -224 11960 -197 11985
rect -157 11960 -154 11985
rect -154 11960 -123 11985
rect -305 11951 -271 11960
rect -231 11951 -197 11960
rect -157 11951 -123 11960
rect -818 11892 -784 11925
rect -305 11892 -294 11913
rect -294 11892 -271 11913
rect -231 11892 -224 11913
rect -224 11892 -197 11913
rect -157 11892 -154 11913
rect -154 11892 -123 11913
rect -818 11891 -784 11892
rect -305 11879 -271 11892
rect -231 11879 -197 11892
rect -157 11879 -123 11892
rect -818 11824 -784 11853
rect -305 11824 -294 11841
rect -294 11824 -271 11841
rect -231 11824 -224 11841
rect -224 11824 -197 11841
rect -157 11824 -154 11841
rect -154 11824 -123 11841
rect -818 11819 -784 11824
rect -305 11807 -271 11824
rect -231 11807 -197 11824
rect -157 11807 -123 11824
rect -818 11756 -784 11781
rect -305 11756 -294 11769
rect -294 11756 -271 11769
rect -231 11756 -224 11769
rect -224 11756 -197 11769
rect -157 11756 -154 11769
rect -154 11756 -123 11769
rect -818 11747 -784 11756
rect -305 11735 -271 11756
rect -231 11735 -197 11756
rect -157 11735 -123 11756
rect -818 11688 -784 11709
rect -305 11688 -294 11697
rect -294 11688 -271 11697
rect -231 11688 -224 11697
rect -224 11688 -197 11697
rect -157 11688 -154 11697
rect -154 11688 -123 11697
rect -818 11675 -784 11688
rect -305 11663 -271 11688
rect -231 11663 -197 11688
rect -157 11663 -123 11688
rect -818 11620 -784 11637
rect -305 11620 -294 11625
rect -294 11620 -271 11625
rect -231 11620 -224 11625
rect -224 11620 -197 11625
rect -157 11620 -154 11625
rect -154 11620 -123 11625
rect -818 11603 -784 11620
rect -305 11591 -271 11620
rect -231 11591 -197 11620
rect -157 11591 -123 11620
rect -818 11552 -784 11565
rect -305 11552 -294 11553
rect -294 11552 -271 11553
rect -231 11552 -224 11553
rect -224 11552 -197 11553
rect -157 11552 -154 11553
rect -154 11552 -123 11553
rect -818 11531 -784 11552
rect -305 11519 -271 11552
rect -231 11519 -197 11552
rect -157 11519 -123 11552
rect -818 11484 -784 11493
rect -818 11459 -784 11484
rect -305 11450 -271 11481
rect -231 11450 -197 11481
rect -157 11450 -123 11481
rect -818 11416 -784 11421
rect -305 11447 -294 11450
rect -294 11447 -271 11450
rect -231 11447 -224 11450
rect -224 11447 -197 11450
rect -157 11447 -154 11450
rect -154 11447 -123 11450
rect -818 11387 -784 11416
rect -305 11382 -271 11409
rect -231 11382 -197 11409
rect -157 11382 -123 11409
rect -818 11348 -784 11349
rect -305 11375 -294 11382
rect -294 11375 -271 11382
rect -231 11375 -224 11382
rect -224 11375 -197 11382
rect -157 11375 -154 11382
rect -154 11375 -123 11382
rect -818 11315 -784 11348
rect -305 11314 -271 11337
rect -231 11314 -197 11337
rect -157 11314 -123 11337
rect -305 11303 -294 11314
rect -294 11303 -271 11314
rect -231 11303 -224 11314
rect -224 11303 -197 11314
rect -157 11303 -154 11314
rect -154 11303 -123 11314
rect -818 11246 -784 11277
rect -305 11246 -271 11265
rect -231 11246 -197 11265
rect -157 11246 -123 11265
rect -818 11243 -784 11246
rect -305 11231 -294 11246
rect -294 11231 -271 11246
rect -231 11231 -224 11246
rect -224 11231 -197 11246
rect -157 11231 -154 11246
rect -154 11231 -123 11246
rect -818 11178 -784 11205
rect -305 11178 -271 11193
rect -231 11178 -197 11193
rect -157 11178 -123 11193
rect -818 11171 -784 11178
rect -305 11159 -294 11178
rect -294 11159 -271 11178
rect -231 11159 -224 11178
rect -224 11159 -197 11178
rect -157 11159 -154 11178
rect -154 11159 -123 11178
rect -818 11110 -784 11133
rect -305 11110 -271 11121
rect -231 11110 -197 11121
rect -157 11110 -123 11121
rect -818 11099 -784 11110
rect -305 11087 -294 11110
rect -294 11087 -271 11110
rect -231 11087 -224 11110
rect -224 11087 -197 11110
rect -157 11087 -154 11110
rect -154 11087 -123 11110
rect -818 11042 -784 11061
rect -305 11042 -271 11049
rect -231 11042 -197 11049
rect -157 11042 -123 11049
rect -818 11027 -784 11042
rect -305 11015 -294 11042
rect -294 11015 -271 11042
rect -231 11015 -224 11042
rect -224 11015 -197 11042
rect -157 11015 -154 11042
rect -154 11015 -123 11042
rect -818 10974 -784 10989
rect -305 10974 -271 10977
rect -231 10974 -197 10977
rect -157 10974 -123 10977
rect -818 10955 -784 10974
rect -305 10943 -294 10974
rect -294 10943 -271 10974
rect -231 10943 -224 10974
rect -224 10943 -197 10974
rect -157 10943 -154 10974
rect -154 10943 -123 10974
rect -818 10906 -784 10917
rect -818 10883 -784 10906
rect -305 10872 -294 10905
rect -294 10872 -271 10905
rect -231 10872 -224 10905
rect -224 10872 -197 10905
rect -157 10872 -154 10905
rect -154 10872 -123 10905
rect -305 10871 -271 10872
rect -231 10871 -197 10872
rect -157 10871 -123 10872
rect -818 10838 -784 10845
rect -818 10811 -784 10838
rect -305 10804 -294 10833
rect -294 10804 -271 10833
rect -231 10804 -224 10833
rect -224 10804 -197 10833
rect -157 10804 -154 10833
rect -154 10804 -123 10833
rect -305 10799 -271 10804
rect -231 10799 -197 10804
rect -157 10799 -123 10804
rect -818 10770 -784 10773
rect -818 10739 -784 10770
rect -305 10736 -294 10761
rect -294 10736 -271 10761
rect -231 10736 -224 10761
rect -224 10736 -197 10761
rect -157 10736 -154 10761
rect -154 10736 -123 10761
rect -305 10727 -271 10736
rect -231 10727 -197 10736
rect -157 10727 -123 10736
rect -818 10668 -784 10701
rect -305 10668 -294 10689
rect -294 10668 -271 10689
rect -231 10668 -224 10689
rect -224 10668 -197 10689
rect -157 10668 -154 10689
rect -154 10668 -123 10689
rect -818 10667 -784 10668
rect -305 10655 -271 10668
rect -231 10655 -197 10668
rect -157 10655 -123 10668
rect -818 10600 -784 10629
rect -305 10600 -294 10617
rect -294 10600 -271 10617
rect -231 10600 -224 10617
rect -224 10600 -197 10617
rect -157 10600 -154 10617
rect -154 10600 -123 10617
rect -818 10595 -784 10600
rect -305 10583 -271 10600
rect -231 10583 -197 10600
rect -157 10583 -123 10600
rect -818 10532 -784 10557
rect -305 10532 -294 10545
rect -294 10532 -271 10545
rect -231 10532 -224 10545
rect -224 10532 -197 10545
rect -157 10532 -154 10545
rect -154 10532 -123 10545
rect -818 10523 -784 10532
rect -305 10511 -271 10532
rect -231 10511 -197 10532
rect -157 10511 -123 10532
rect -818 10464 -784 10485
rect -305 10464 -294 10473
rect -294 10464 -271 10473
rect -231 10464 -224 10473
rect -224 10464 -197 10473
rect -157 10464 -154 10473
rect -154 10464 -123 10473
rect -818 10451 -784 10464
rect -305 10439 -271 10464
rect -231 10439 -197 10464
rect -157 10439 -123 10464
rect -818 10396 -784 10413
rect -305 10396 -294 10401
rect -294 10396 -271 10401
rect -231 10396 -224 10401
rect -224 10396 -197 10401
rect -157 10396 -154 10401
rect -154 10396 -123 10401
rect -818 10379 -784 10396
rect -305 10367 -271 10396
rect -231 10367 -197 10396
rect -157 10367 -123 10396
rect -818 10328 -784 10341
rect -305 10328 -294 10329
rect -294 10328 -271 10329
rect -231 10328 -224 10329
rect -224 10328 -197 10329
rect -157 10328 -154 10329
rect -154 10328 -123 10329
rect -818 10307 -784 10328
rect -305 10295 -271 10328
rect -231 10295 -197 10328
rect -157 10295 -123 10328
rect -818 10260 -784 10269
rect -818 10235 -784 10260
rect -305 10226 -271 10257
rect -231 10226 -197 10257
rect -157 10226 -123 10257
rect -818 10192 -784 10197
rect -305 10223 -294 10226
rect -294 10223 -271 10226
rect -231 10223 -224 10226
rect -224 10223 -197 10226
rect -157 10223 -154 10226
rect -154 10223 -123 10226
rect -818 10163 -784 10192
rect -305 10158 -271 10185
rect -231 10158 -197 10185
rect -157 10158 -123 10185
rect -818 10124 -784 10125
rect -305 10151 -294 10158
rect -294 10151 -271 10158
rect -231 10151 -224 10158
rect -224 10151 -197 10158
rect -157 10151 -154 10158
rect -154 10151 -123 10158
rect -818 10091 -784 10124
rect -305 10090 -271 10113
rect -231 10090 -197 10113
rect -157 10090 -123 10113
rect -305 10079 -294 10090
rect -294 10079 -271 10090
rect -231 10079 -224 10090
rect -224 10079 -197 10090
rect -157 10079 -154 10090
rect -154 10079 -123 10090
rect -818 10022 -784 10053
rect -305 10022 -271 10041
rect -231 10022 -197 10041
rect -157 10022 -123 10041
rect -818 10019 -784 10022
rect -305 10007 -294 10022
rect -294 10007 -271 10022
rect -231 10007 -224 10022
rect -224 10007 -197 10022
rect -157 10007 -154 10022
rect -154 10007 -123 10022
rect -818 9954 -784 9981
rect -305 9954 -271 9969
rect -231 9954 -197 9969
rect -157 9954 -123 9969
rect -818 9947 -784 9954
rect -305 9935 -294 9954
rect -294 9935 -271 9954
rect -231 9935 -224 9954
rect -224 9935 -197 9954
rect -157 9935 -154 9954
rect -154 9935 -123 9954
rect -818 9886 -784 9909
rect -305 9886 -271 9897
rect -231 9886 -197 9897
rect -157 9886 -123 9897
rect -818 9875 -784 9886
rect -305 9863 -294 9886
rect -294 9863 -271 9886
rect -231 9863 -224 9886
rect -224 9863 -197 9886
rect -157 9863 -154 9886
rect -154 9863 -123 9886
rect -818 9818 -784 9837
rect -305 9818 -271 9825
rect -231 9818 -197 9825
rect -157 9818 -123 9825
rect -818 9803 -784 9818
rect -305 9791 -294 9818
rect -294 9791 -271 9818
rect -231 9791 -224 9818
rect -224 9791 -197 9818
rect -157 9791 -154 9818
rect -154 9791 -123 9818
rect -818 9750 -784 9765
rect -305 9750 -271 9753
rect -231 9750 -197 9753
rect -157 9750 -123 9753
rect -818 9731 -784 9750
rect -305 9719 -294 9750
rect -294 9719 -271 9750
rect -231 9719 -224 9750
rect -224 9719 -197 9750
rect -157 9719 -154 9750
rect -154 9719 -123 9750
rect -818 9682 -784 9693
rect -818 9659 -784 9682
rect -305 9648 -294 9681
rect -294 9648 -271 9681
rect -231 9648 -224 9681
rect -224 9648 -197 9681
rect -157 9648 -154 9681
rect -154 9648 -123 9681
rect -305 9647 -271 9648
rect -231 9647 -197 9648
rect -157 9647 -123 9648
rect -818 9614 -784 9621
rect -818 9587 -784 9614
rect -305 9580 -294 9609
rect -294 9580 -271 9609
rect -231 9580 -224 9609
rect -224 9580 -197 9609
rect -157 9580 -154 9609
rect -154 9580 -123 9609
rect -305 9575 -271 9580
rect -231 9575 -197 9580
rect -157 9575 -123 9580
rect -818 9546 -784 9549
rect -818 9515 -784 9546
rect -305 9512 -294 9537
rect -294 9512 -271 9537
rect -231 9512 -224 9537
rect -224 9512 -197 9537
rect -157 9512 -154 9537
rect -154 9512 -123 9537
rect -305 9503 -271 9512
rect -231 9503 -197 9512
rect -157 9503 -123 9512
rect -818 9444 -784 9477
rect -305 9444 -294 9465
rect -294 9444 -271 9465
rect -231 9444 -224 9465
rect -224 9444 -197 9465
rect -157 9444 -154 9465
rect -154 9444 -123 9465
rect -818 9443 -784 9444
rect -305 9431 -271 9444
rect -231 9431 -197 9444
rect -157 9431 -123 9444
rect -818 9376 -784 9405
rect -305 9376 -294 9393
rect -294 9376 -271 9393
rect -231 9376 -224 9393
rect -224 9376 -197 9393
rect -157 9376 -154 9393
rect -154 9376 -123 9393
rect -818 9371 -784 9376
rect -305 9359 -271 9376
rect -231 9359 -197 9376
rect -157 9359 -123 9376
rect -818 9308 -784 9333
rect -305 9308 -294 9321
rect -294 9308 -271 9321
rect -231 9308 -224 9321
rect -224 9308 -197 9321
rect -157 9308 -154 9321
rect -154 9308 -123 9321
rect -818 9299 -784 9308
rect -305 9287 -271 9308
rect -231 9287 -197 9308
rect -157 9287 -123 9308
rect -818 9240 -784 9261
rect -305 9240 -294 9249
rect -294 9240 -271 9249
rect -231 9240 -224 9249
rect -224 9240 -197 9249
rect -157 9240 -154 9249
rect -154 9240 -123 9249
rect -818 9227 -784 9240
rect -305 9215 -271 9240
rect -231 9215 -197 9240
rect -157 9215 -123 9240
rect -818 9172 -784 9189
rect -305 9172 -294 9177
rect -294 9172 -271 9177
rect -231 9172 -224 9177
rect -224 9172 -197 9177
rect -157 9172 -154 9177
rect -154 9172 -123 9177
rect -818 9155 -784 9172
rect -305 9143 -271 9172
rect -231 9143 -197 9172
rect -157 9143 -123 9172
rect -818 9104 -784 9117
rect -305 9104 -294 9105
rect -294 9104 -271 9105
rect -231 9104 -224 9105
rect -224 9104 -197 9105
rect -157 9104 -154 9105
rect -154 9104 -123 9105
rect -818 9083 -784 9104
rect -305 9071 -271 9104
rect -231 9071 -197 9104
rect -157 9071 -123 9104
rect -818 9036 -784 9045
rect -818 9011 -784 9036
rect -305 9002 -271 9033
rect -231 9002 -197 9033
rect -157 9002 -123 9033
rect -818 8968 -784 8973
rect -305 8999 -294 9002
rect -294 8999 -271 9002
rect -231 8999 -224 9002
rect -224 8999 -197 9002
rect -157 8999 -154 9002
rect -154 8999 -123 9002
rect -818 8939 -784 8968
rect -305 8934 -271 8961
rect -231 8934 -197 8961
rect -157 8934 -123 8961
rect -818 8900 -784 8901
rect -305 8927 -294 8934
rect -294 8927 -271 8934
rect -231 8927 -224 8934
rect -224 8927 -197 8934
rect -157 8927 -154 8934
rect -154 8927 -123 8934
rect -818 8867 -784 8900
rect -305 8866 -271 8889
rect -231 8866 -197 8889
rect -157 8866 -123 8889
rect -305 8855 -294 8866
rect -294 8855 -271 8866
rect -231 8855 -224 8866
rect -224 8855 -197 8866
rect -157 8855 -154 8866
rect -154 8855 -123 8866
rect -818 8798 -784 8829
rect -305 8798 -271 8817
rect -231 8798 -197 8817
rect -157 8798 -123 8817
rect -818 8795 -784 8798
rect -305 8783 -294 8798
rect -294 8783 -271 8798
rect -231 8783 -224 8798
rect -224 8783 -197 8798
rect -157 8783 -154 8798
rect -154 8783 -123 8798
rect -818 8730 -784 8757
rect -305 8730 -271 8745
rect -231 8730 -197 8745
rect -157 8730 -123 8745
rect -818 8723 -784 8730
rect -305 8711 -294 8730
rect -294 8711 -271 8730
rect -231 8711 -224 8730
rect -224 8711 -197 8730
rect -157 8711 -154 8730
rect -154 8711 -123 8730
rect -818 8662 -784 8685
rect -305 8662 -271 8673
rect -231 8662 -197 8673
rect -157 8662 -123 8673
rect -818 8651 -784 8662
rect -305 8639 -294 8662
rect -294 8639 -271 8662
rect -231 8639 -224 8662
rect -224 8639 -197 8662
rect -157 8639 -154 8662
rect -154 8639 -123 8662
rect -818 8594 -784 8613
rect -305 8594 -271 8601
rect -231 8594 -197 8601
rect -157 8594 -123 8601
rect -818 8579 -784 8594
rect -305 8567 -294 8594
rect -294 8567 -271 8594
rect -231 8567 -224 8594
rect -224 8567 -197 8594
rect -157 8567 -154 8594
rect -154 8567 -123 8594
rect -818 8526 -784 8541
rect -305 8526 -271 8529
rect -231 8526 -197 8529
rect -157 8526 -123 8529
rect -818 8507 -784 8526
rect -305 8495 -294 8526
rect -294 8495 -271 8526
rect -231 8495 -224 8526
rect -224 8495 -197 8526
rect -157 8495 -154 8526
rect -154 8495 -123 8526
rect -818 8458 -784 8469
rect -818 8435 -784 8458
rect -305 8424 -294 8457
rect -294 8424 -271 8457
rect -231 8424 -224 8457
rect -224 8424 -197 8457
rect -157 8424 -154 8457
rect -154 8424 -123 8457
rect -305 8423 -271 8424
rect -231 8423 -197 8424
rect -157 8423 -123 8424
rect -818 8390 -784 8397
rect -818 8363 -784 8390
rect -305 8356 -294 8385
rect -294 8356 -271 8385
rect -231 8356 -224 8385
rect -224 8356 -197 8385
rect -157 8356 -154 8385
rect -154 8356 -123 8385
rect -305 8351 -271 8356
rect -231 8351 -197 8356
rect -157 8351 -123 8356
rect -818 8322 -784 8325
rect -818 8291 -784 8322
rect -305 8288 -294 8313
rect -294 8288 -271 8313
rect -231 8288 -224 8313
rect -224 8288 -197 8313
rect -157 8288 -154 8313
rect -154 8288 -123 8313
rect -305 8279 -271 8288
rect -231 8279 -197 8288
rect -157 8279 -123 8288
rect -818 8220 -784 8253
rect -305 8220 -294 8241
rect -294 8220 -271 8241
rect -231 8220 -224 8241
rect -224 8220 -197 8241
rect -157 8220 -154 8241
rect -154 8220 -123 8241
rect -818 8219 -784 8220
rect -305 8207 -271 8220
rect -231 8207 -197 8220
rect -157 8207 -123 8220
rect -818 8152 -784 8181
rect -305 8152 -294 8168
rect -294 8152 -271 8168
rect -231 8152 -224 8168
rect -224 8152 -197 8168
rect -157 8152 -154 8168
rect -154 8152 -123 8168
rect -818 8147 -784 8152
rect -305 8134 -271 8152
rect -231 8134 -197 8152
rect -157 8134 -123 8152
rect -818 8084 -784 8109
rect -305 8084 -294 8095
rect -294 8084 -271 8095
rect -231 8084 -224 8095
rect -224 8084 -197 8095
rect -157 8084 -154 8095
rect -154 8084 -123 8095
rect -818 8075 -784 8084
rect -305 8061 -271 8084
rect -231 8061 -197 8084
rect -157 8061 -123 8084
rect -818 8016 -784 8037
rect -305 8016 -294 8022
rect -294 8016 -271 8022
rect -231 8016 -224 8022
rect -224 8016 -197 8022
rect -157 8016 -154 8022
rect -154 8016 -123 8022
rect -818 8003 -784 8016
rect -305 7988 -271 8016
rect -231 7988 -197 8016
rect -157 7988 -123 8016
rect -818 7948 -784 7965
rect -305 7948 -294 7949
rect -294 7948 -271 7949
rect -231 7948 -224 7949
rect -224 7948 -197 7949
rect -157 7948 -154 7949
rect -154 7948 -123 7949
rect -818 7931 -784 7948
rect -305 7915 -271 7948
rect -231 7915 -197 7948
rect -157 7915 -123 7948
rect -818 7880 -784 7893
rect -818 7859 -784 7880
rect -305 7846 -271 7876
rect -231 7846 -197 7876
rect -157 7846 -123 7876
rect -818 7812 -784 7821
rect -305 7842 -294 7846
rect -294 7842 -271 7846
rect -231 7842 -224 7846
rect -224 7842 -197 7846
rect -157 7842 -154 7846
rect -154 7842 -123 7846
rect -818 7787 -784 7812
rect -305 7778 -271 7803
rect -231 7778 -197 7803
rect -157 7778 -123 7803
rect -818 7744 -784 7749
rect -305 7769 -294 7778
rect -294 7769 -271 7778
rect -231 7769 -224 7778
rect -224 7769 -197 7778
rect -157 7769 -154 7778
rect -154 7769 -123 7778
rect -818 7715 -784 7744
rect -305 7710 -271 7730
rect -231 7710 -197 7730
rect -157 7710 -123 7730
rect -818 7676 -784 7677
rect -305 7696 -294 7710
rect -294 7696 -271 7710
rect -231 7696 -224 7710
rect -224 7696 -197 7710
rect -157 7696 -154 7710
rect -154 7696 -123 7710
rect -818 7643 -784 7676
rect -305 7642 -271 7657
rect -231 7642 -197 7657
rect -157 7642 -123 7657
rect -305 7623 -294 7642
rect -294 7623 -271 7642
rect -231 7623 -224 7642
rect -224 7623 -197 7642
rect -157 7623 -154 7642
rect -154 7623 -123 7642
rect -818 7574 -784 7605
rect -305 7574 -271 7584
rect -231 7574 -197 7584
rect -157 7574 -123 7584
rect -818 7571 -784 7574
rect -305 7550 -294 7574
rect -294 7550 -271 7574
rect -231 7550 -224 7574
rect -224 7550 -197 7574
rect -157 7550 -154 7574
rect -154 7550 -123 7574
rect -818 7506 -784 7533
rect -305 7506 -271 7511
rect -231 7506 -197 7511
rect -157 7506 -123 7511
rect -818 7499 -784 7506
rect -305 7477 -294 7506
rect -294 7477 -271 7506
rect -231 7477 -224 7506
rect -224 7477 -197 7506
rect -157 7477 -154 7506
rect -154 7477 -123 7506
rect -818 7438 -784 7461
rect -818 7427 -784 7438
rect -305 7404 -294 7438
rect -294 7404 -271 7438
rect -231 7404 -224 7438
rect -224 7404 -197 7438
rect -157 7404 -154 7438
rect -154 7404 -123 7438
rect -818 7370 -784 7389
rect -818 7355 -784 7370
rect -305 7336 -294 7365
rect -294 7336 -271 7365
rect -231 7336 -224 7365
rect -224 7336 -197 7365
rect -157 7336 -154 7365
rect -154 7336 -123 7365
rect -305 7331 -271 7336
rect -231 7331 -197 7336
rect -157 7331 -123 7336
rect -818 7302 -784 7317
rect -818 7283 -784 7302
rect -305 7268 -294 7292
rect -294 7268 -271 7292
rect -231 7268 -224 7292
rect -224 7268 -197 7292
rect -157 7268 -154 7292
rect -154 7268 -123 7292
rect -305 7258 -271 7268
rect -231 7258 -197 7268
rect -157 7258 -123 7268
rect -818 7234 -784 7245
rect -818 7211 -784 7234
rect -305 7200 -294 7219
rect -294 7200 -271 7219
rect -231 7200 -224 7219
rect -224 7200 -197 7219
rect -157 7200 -154 7219
rect -154 7200 -123 7219
rect -305 7185 -271 7200
rect -231 7185 -197 7200
rect -157 7185 -123 7200
rect -818 7166 -784 7173
rect -818 7139 -784 7166
rect -305 7132 -294 7146
rect -294 7132 -271 7146
rect -231 7132 -224 7146
rect -224 7132 -197 7146
rect -157 7132 -154 7146
rect -154 7132 -123 7146
rect -305 7112 -271 7132
rect -231 7112 -197 7132
rect -157 7112 -123 7132
rect -818 7098 -784 7101
rect -818 7067 -784 7098
rect -305 7064 -294 7073
rect -294 7064 -271 7073
rect -231 7064 -224 7073
rect -224 7064 -197 7073
rect -157 7064 -154 7073
rect -154 7064 -123 7073
rect -305 7039 -271 7064
rect -231 7039 -197 7064
rect -157 7039 -123 7064
rect -818 6996 -784 7029
rect -305 6996 -294 7000
rect -294 6996 -271 7000
rect -231 6996 -224 7000
rect -224 6996 -197 7000
rect -157 6996 -154 7000
rect -154 6996 -123 7000
rect -818 6995 -784 6996
rect -305 6966 -271 6996
rect -231 6966 -197 6996
rect -157 6966 -123 6996
rect -818 6928 -784 6957
rect -818 6923 -784 6928
rect -305 6894 -271 6927
rect -231 6894 -197 6927
rect -157 6894 -123 6927
rect -818 6860 -784 6885
rect -305 6893 -294 6894
rect -294 6893 -271 6894
rect -231 6893 -224 6894
rect -224 6893 -197 6894
rect -157 6893 -154 6894
rect -154 6893 -123 6894
rect -818 6851 -784 6860
rect -305 6826 -271 6854
rect -231 6826 -197 6854
rect -157 6826 -123 6854
rect -818 6792 -784 6813
rect -305 6820 -294 6826
rect -294 6820 -271 6826
rect -231 6820 -224 6826
rect -224 6820 -197 6826
rect -157 6820 -154 6826
rect -154 6820 -123 6826
rect -818 6779 -784 6792
rect -305 6758 -271 6781
rect -231 6758 -197 6781
rect -157 6758 -123 6781
rect -818 6724 -784 6741
rect -305 6747 -294 6758
rect -294 6747 -271 6758
rect -231 6747 -224 6758
rect -224 6747 -197 6758
rect -157 6747 -154 6758
rect -154 6747 -123 6758
rect -818 6707 -784 6724
rect -305 6690 -271 6708
rect -231 6690 -197 6708
rect -157 6690 -123 6708
rect -818 6656 -784 6669
rect -305 6674 -294 6690
rect -294 6674 -271 6690
rect -231 6674 -224 6690
rect -224 6674 -197 6690
rect -157 6674 -154 6690
rect -154 6674 -123 6690
rect -818 6635 -784 6656
rect -305 6622 -271 6635
rect -231 6622 -197 6635
rect -157 6622 -123 6635
rect -818 6588 -784 6597
rect -305 6601 -294 6622
rect -294 6601 -271 6622
rect -231 6601 -224 6622
rect -224 6601 -197 6622
rect -157 6601 -154 6622
rect -154 6601 -123 6622
rect -818 6563 -784 6588
rect -305 6554 -271 6562
rect -231 6554 -197 6562
rect -157 6554 -123 6562
rect -818 6520 -784 6525
rect -305 6528 -294 6554
rect -294 6528 -271 6554
rect -231 6528 -224 6554
rect -224 6528 -197 6554
rect -157 6528 -154 6554
rect -154 6528 -123 6554
rect -818 6491 -784 6520
rect -305 6486 -271 6489
rect -231 6486 -197 6489
rect -157 6486 -123 6489
rect -818 6452 -784 6453
rect -305 6455 -294 6486
rect -294 6455 -271 6486
rect -231 6455 -224 6486
rect -224 6455 -197 6486
rect -157 6455 -154 6486
rect -154 6455 -123 6486
rect -818 6419 -784 6452
rect -305 6384 -294 6416
rect -294 6384 -271 6416
rect -231 6384 -224 6416
rect -224 6384 -197 6416
rect -157 6384 -154 6416
rect -154 6384 -123 6416
rect -305 6382 -271 6384
rect -231 6382 -197 6384
rect -157 6382 -123 6384
rect -818 6350 -784 6381
rect -818 6347 -784 6350
rect -305 6316 -294 6343
rect -294 6316 -271 6343
rect -231 6316 -224 6343
rect -224 6316 -197 6343
rect -157 6316 -154 6343
rect -154 6316 -123 6343
rect -305 6309 -271 6316
rect -231 6309 -197 6316
rect -157 6309 -123 6316
rect -818 6282 -784 6309
rect -818 6275 -784 6282
rect -305 6248 -294 6270
rect -294 6248 -271 6270
rect -231 6248 -224 6270
rect -224 6248 -197 6270
rect -157 6248 -154 6270
rect -154 6248 -123 6270
rect -818 6214 -784 6237
rect -305 6236 -271 6248
rect -231 6236 -197 6248
rect -157 6236 -123 6248
rect -818 6203 -784 6214
rect -305 6180 -294 6197
rect -294 6180 -271 6197
rect -231 6180 -224 6197
rect -224 6180 -197 6197
rect -157 6180 -154 6197
rect -154 6180 -123 6197
rect -818 6146 -784 6165
rect -305 6163 -271 6180
rect -231 6163 -197 6180
rect -157 6163 -123 6180
rect -818 6131 -784 6146
rect -305 6112 -294 6124
rect -294 6112 -271 6124
rect -231 6112 -224 6124
rect -224 6112 -197 6124
rect -157 6112 -154 6124
rect -154 6112 -123 6124
rect -818 6078 -784 6093
rect -305 6090 -271 6112
rect -231 6090 -197 6112
rect -157 6090 -123 6112
rect -818 6059 -784 6078
rect -305 6044 -294 6051
rect -294 6044 -271 6051
rect -231 6044 -224 6051
rect -224 6044 -197 6051
rect -157 6044 -154 6051
rect -154 6044 -123 6051
rect -818 6010 -784 6021
rect -305 6017 -271 6044
rect -231 6017 -197 6044
rect -157 6017 -123 6044
rect -818 5987 -784 6010
rect -305 5976 -294 5978
rect -294 5976 -271 5978
rect -231 5976 -224 5978
rect -224 5976 -197 5978
rect -157 5976 -154 5978
rect -154 5976 -123 5978
rect -818 5942 -784 5949
rect -305 5944 -271 5976
rect -231 5944 -197 5976
rect -157 5944 -123 5976
rect -818 5915 -784 5942
rect -818 5874 -784 5877
rect -305 5874 -271 5905
rect -231 5874 -197 5905
rect -157 5874 -123 5905
rect -818 5843 -784 5874
rect -305 5871 -294 5874
rect -294 5871 -271 5874
rect -231 5871 -224 5874
rect -224 5871 -197 5874
rect -157 5871 -154 5874
rect -154 5871 -123 5874
rect -305 5806 -271 5832
rect -231 5806 -197 5832
rect -157 5806 -123 5832
rect -818 5772 -784 5805
rect -305 5798 -294 5806
rect -294 5798 -271 5806
rect -231 5798 -224 5806
rect -224 5798 -197 5806
rect -157 5798 -154 5806
rect -154 5798 -123 5806
rect -818 5771 -784 5772
rect -305 5738 -271 5759
rect -231 5738 -197 5759
rect -157 5738 -123 5759
rect -818 5704 -784 5733
rect -305 5725 -294 5738
rect -294 5725 -271 5738
rect -231 5725 -224 5738
rect -224 5725 -197 5738
rect -157 5725 -154 5738
rect -154 5725 -123 5738
rect -818 5699 -784 5704
rect -305 5670 -271 5686
rect -231 5670 -197 5686
rect -157 5670 -123 5686
rect -818 5636 -784 5661
rect -305 5652 -294 5670
rect -294 5652 -271 5670
rect -231 5652 -224 5670
rect -224 5652 -197 5670
rect -157 5652 -154 5670
rect -154 5652 -123 5670
rect -818 5627 -784 5636
rect -305 5602 -271 5613
rect -231 5602 -197 5613
rect -157 5602 -123 5613
rect -818 5568 -784 5589
rect -305 5579 -294 5602
rect -294 5579 -271 5602
rect -231 5579 -224 5602
rect -224 5579 -197 5602
rect -157 5579 -154 5602
rect -154 5579 -123 5602
rect -818 5555 -784 5568
rect -305 5534 -271 5540
rect -231 5534 -197 5540
rect -157 5534 -123 5540
rect -818 5500 -784 5517
rect -305 5506 -294 5534
rect -294 5506 -271 5534
rect -231 5506 -224 5534
rect -224 5506 -197 5534
rect -157 5506 -154 5534
rect -154 5506 -123 5534
rect -818 5483 -784 5500
rect -305 5466 -271 5467
rect -231 5466 -197 5467
rect -157 5466 -123 5467
rect -818 5432 -784 5445
rect -305 5433 -294 5466
rect -294 5433 -271 5466
rect -231 5433 -224 5466
rect -224 5433 -197 5466
rect -157 5433 -154 5466
rect -154 5433 -123 5466
rect -818 5411 -784 5432
rect -818 5364 -784 5373
rect -305 5364 -294 5394
rect -294 5364 -271 5394
rect -231 5364 -224 5394
rect -224 5364 -197 5394
rect -157 5364 -154 5394
rect -154 5364 -123 5394
rect -818 5339 -784 5364
rect -305 5360 -271 5364
rect -231 5360 -197 5364
rect -157 5360 -123 5364
rect -818 5296 -784 5301
rect -305 5296 -294 5321
rect -294 5296 -271 5321
rect -231 5296 -224 5321
rect -224 5296 -197 5321
rect -157 5296 -154 5321
rect -154 5296 -123 5321
rect -818 5267 -784 5296
rect -305 5287 -271 5296
rect -231 5287 -197 5296
rect -157 5287 -123 5296
rect -818 5228 -784 5229
rect -305 5228 -294 5248
rect -294 5228 -271 5248
rect -231 5228 -224 5248
rect -224 5228 -197 5248
rect -157 5228 -154 5248
rect -154 5228 -123 5248
rect -818 5195 -784 5228
rect -305 5214 -271 5228
rect -231 5214 -197 5228
rect -157 5214 -123 5228
rect -305 5160 -294 5175
rect -294 5160 -271 5175
rect -231 5160 -224 5175
rect -224 5160 -197 5175
rect -157 5160 -154 5175
rect -154 5160 -123 5175
rect -818 5126 -784 5157
rect -305 5141 -271 5160
rect -231 5141 -197 5160
rect -157 5141 -123 5160
rect -818 5123 -784 5126
rect -305 5092 -294 5102
rect -294 5092 -271 5102
rect -231 5092 -224 5102
rect -224 5092 -197 5102
rect -157 5092 -154 5102
rect -154 5092 -123 5102
rect -818 5058 -784 5085
rect -305 5068 -271 5092
rect -231 5068 -197 5092
rect -157 5068 -123 5092
rect -818 5051 -784 5058
rect -305 5024 -294 5029
rect -294 5024 -271 5029
rect -231 5024 -224 5029
rect -224 5024 -197 5029
rect -157 5024 -154 5029
rect -154 5024 -123 5029
rect -818 4990 -784 5013
rect -305 4995 -271 5024
rect -231 4995 -197 5024
rect -157 4995 -123 5024
rect -818 4979 -784 4990
rect 28 4976 62 5010
rect -62 4956 -48 4974
rect -48 4956 -28 4974
rect -818 4922 -784 4941
rect -305 4922 -271 4956
rect -231 4922 -197 4956
rect -157 4922 -123 4956
rect -62 4940 -28 4956
rect 106 4976 140 5010
rect 184 4976 218 5010
rect 262 4976 296 5010
rect 340 4976 374 5010
rect 418 4976 452 5010
rect 496 4976 530 5010
rect 574 4976 608 5010
rect 652 4976 686 5010
rect 730 4976 764 5010
rect 808 4976 842 5010
rect -818 4907 -784 4922
rect -62 4888 -48 4901
rect -48 4888 -28 4901
rect -818 4854 -784 4869
rect -305 4854 -271 4883
rect -231 4854 -197 4883
rect -157 4854 -123 4883
rect -62 4867 -28 4888
rect -818 4835 -784 4854
rect -305 4849 -294 4854
rect -294 4849 -271 4854
rect -231 4849 -224 4854
rect -224 4849 -197 4854
rect -157 4849 -154 4854
rect -154 4849 -123 4854
rect -62 4820 -48 4828
rect -48 4820 -28 4828
rect -818 4786 -784 4797
rect -305 4786 -271 4810
rect -231 4786 -197 4810
rect -157 4786 -123 4810
rect -62 4794 -28 4820
rect -818 4763 -784 4786
rect -305 4776 -294 4786
rect -294 4776 -271 4786
rect -231 4776 -224 4786
rect -224 4776 -197 4786
rect -157 4776 -154 4786
rect -154 4776 -123 4786
rect -62 4752 -48 4755
rect -48 4752 -28 4755
rect -818 4718 -784 4725
rect -305 4718 -271 4737
rect -231 4718 -197 4737
rect -157 4718 -123 4737
rect -62 4721 -28 4752
rect -818 4691 -784 4718
rect -305 4703 -294 4718
rect -294 4703 -271 4718
rect -231 4703 -224 4718
rect -224 4703 -197 4718
rect -157 4703 -154 4718
rect -154 4703 -123 4718
rect -818 4650 -784 4653
rect -305 4650 -271 4664
rect -231 4650 -197 4664
rect -157 4650 -123 4664
rect -62 4650 -28 4682
rect -818 4619 -784 4650
rect -305 4630 -294 4650
rect -294 4630 -271 4650
rect -231 4630 -224 4650
rect -224 4630 -197 4650
rect -157 4630 -154 4650
rect -154 4630 -123 4650
rect -62 4648 -48 4650
rect -48 4648 -28 4650
rect -305 4582 -271 4591
rect -231 4582 -197 4591
rect -157 4582 -123 4591
rect -62 4582 -28 4609
rect -818 4548 -784 4581
rect -305 4557 -294 4582
rect -294 4557 -271 4582
rect -231 4557 -224 4582
rect -224 4557 -197 4582
rect -157 4557 -154 4582
rect -154 4557 -123 4582
rect -62 4575 -48 4582
rect -48 4575 -28 4582
rect -818 4547 -784 4548
rect -305 4514 -271 4518
rect -231 4514 -197 4518
rect -157 4514 -123 4518
rect -62 4514 -28 4536
rect -818 4480 -784 4509
rect -305 4484 -294 4514
rect -294 4484 -271 4514
rect -231 4484 -224 4514
rect -224 4484 -197 4514
rect -157 4484 -154 4514
rect -154 4484 -123 4514
rect -62 4502 -48 4514
rect -48 4502 -28 4514
rect -818 4475 -784 4480
rect -62 4446 -28 4463
rect -818 4412 -784 4437
rect -305 4412 -294 4445
rect -294 4412 -271 4445
rect -231 4412 -224 4445
rect -224 4412 -197 4445
rect -157 4412 -154 4445
rect -154 4412 -123 4445
rect -62 4429 -48 4446
rect -48 4429 -28 4446
rect -818 4403 -784 4412
rect -305 4411 -271 4412
rect -231 4411 -197 4412
rect -157 4411 -123 4412
rect -62 4378 -28 4390
rect -818 4344 -784 4365
rect -305 4344 -294 4372
rect -294 4344 -271 4372
rect -231 4344 -224 4372
rect -224 4344 -197 4372
rect -157 4344 -154 4372
rect -154 4344 -123 4372
rect -62 4356 -48 4378
rect -48 4356 -28 4378
rect -818 4331 -784 4344
rect -305 4338 -271 4344
rect -231 4338 -197 4344
rect -157 4338 -123 4344
rect -62 4310 -28 4317
rect -818 4276 -784 4293
rect -305 4276 -294 4299
rect -294 4276 -271 4299
rect -231 4276 -224 4299
rect -224 4276 -197 4299
rect -157 4276 -154 4299
rect -154 4276 -123 4299
rect -62 4283 -48 4310
rect -48 4283 -28 4310
rect -818 4259 -784 4276
rect -305 4265 -271 4276
rect -231 4265 -197 4276
rect -157 4265 -123 4276
rect -62 4242 -28 4244
rect -818 4208 -784 4221
rect -305 4208 -294 4226
rect -294 4208 -271 4226
rect -231 4208 -224 4226
rect -224 4208 -197 4226
rect -157 4208 -154 4226
rect -154 4208 -123 4226
rect -62 4210 -48 4242
rect -48 4210 -28 4242
rect -818 4187 -784 4208
rect -305 4192 -271 4208
rect -231 4192 -197 4208
rect -157 4192 -123 4208
rect -818 4140 -784 4149
rect -305 4140 -294 4153
rect -294 4140 -271 4153
rect -231 4140 -224 4153
rect -224 4140 -197 4153
rect -157 4140 -154 4153
rect -154 4140 -123 4153
rect -62 4140 -48 4171
rect -48 4140 -28 4171
rect -818 4115 -784 4140
rect -305 4119 -271 4140
rect -231 4119 -197 4140
rect -157 4119 -123 4140
rect -62 4137 -28 4140
rect -818 4072 -784 4077
rect -305 4072 -294 4080
rect -294 4072 -271 4080
rect -231 4072 -224 4080
rect -224 4072 -197 4080
rect -157 4072 -154 4080
rect -154 4072 -123 4080
rect -62 4072 -48 4098
rect -48 4072 -28 4098
rect -818 4043 -784 4072
rect -305 4046 -271 4072
rect -231 4046 -197 4072
rect -157 4046 -123 4072
rect -62 4064 -28 4072
rect -818 4004 -784 4005
rect -305 4004 -294 4007
rect -294 4004 -271 4007
rect -231 4004 -224 4007
rect -224 4004 -197 4007
rect -157 4004 -154 4007
rect -154 4004 -123 4007
rect -62 4004 -48 4026
rect -48 4004 -28 4026
rect -818 3971 -784 4004
rect -305 3973 -271 4004
rect -231 3973 -197 4004
rect -157 3973 -123 4004
rect -62 3992 -28 4004
rect -62 3936 -48 3954
rect -48 3936 -28 3954
rect -818 3902 -784 3933
rect -305 3902 -271 3934
rect -231 3902 -197 3934
rect -157 3902 -123 3934
rect -62 3920 -28 3936
rect -818 3899 -784 3902
rect -305 3900 -294 3902
rect -294 3900 -271 3902
rect -231 3900 -224 3902
rect -224 3900 -197 3902
rect -157 3900 -154 3902
rect -154 3900 -123 3902
rect -62 3868 -48 3882
rect -48 3868 -28 3882
rect -818 3834 -784 3861
rect -305 3834 -271 3861
rect -231 3834 -197 3861
rect -157 3834 -123 3861
rect -62 3848 -28 3868
rect -818 3827 -784 3834
rect -305 3827 -294 3834
rect -294 3827 -271 3834
rect -231 3827 -224 3834
rect -224 3827 -197 3834
rect -157 3827 -154 3834
rect -154 3827 -123 3834
rect -62 3800 -48 3810
rect -48 3800 -28 3810
rect -818 3766 -784 3789
rect -305 3766 -271 3788
rect -231 3766 -197 3788
rect -157 3766 -123 3788
rect -62 3776 -28 3800
rect -818 3755 -784 3766
rect -305 3754 -294 3766
rect -294 3754 -271 3766
rect -231 3754 -224 3766
rect -224 3754 -197 3766
rect -157 3754 -154 3766
rect -154 3754 -123 3766
rect -62 3732 -48 3738
rect -48 3732 -28 3738
rect -818 3698 -784 3717
rect -305 3698 -271 3715
rect -231 3698 -197 3715
rect -157 3698 -123 3715
rect -62 3704 -28 3732
rect -818 3683 -784 3698
rect -305 3681 -294 3698
rect -294 3681 -271 3698
rect -231 3681 -224 3698
rect -224 3681 -197 3698
rect -157 3681 -154 3698
rect -154 3681 -123 3698
rect -62 3664 -48 3666
rect -48 3664 -28 3666
rect -818 3630 -784 3645
rect -305 3630 -271 3642
rect -231 3630 -197 3642
rect -157 3630 -123 3642
rect -62 3632 -28 3664
rect -818 3611 -784 3630
rect -305 3608 -294 3630
rect -294 3608 -271 3630
rect -231 3608 -224 3630
rect -224 3608 -197 3630
rect -157 3608 -154 3630
rect -154 3608 -123 3630
rect -818 3562 -784 3573
rect -305 3562 -271 3569
rect -231 3562 -197 3569
rect -157 3562 -123 3569
rect -62 3562 -28 3594
rect -818 3539 -784 3562
rect -305 3535 -294 3562
rect -294 3535 -271 3562
rect -231 3535 -224 3562
rect -224 3535 -197 3562
rect -157 3535 -154 3562
rect -154 3535 -123 3562
rect -62 3560 -48 3562
rect -48 3560 -28 3562
rect -818 3494 -784 3501
rect -305 3494 -271 3496
rect -231 3494 -197 3496
rect -157 3494 -123 3496
rect -62 3494 -28 3522
rect -818 3467 -784 3494
rect -305 3462 -294 3494
rect -294 3462 -271 3494
rect -231 3462 -224 3494
rect -224 3462 -197 3494
rect -157 3462 -154 3494
rect -154 3462 -123 3494
rect -62 3488 -48 3494
rect -48 3488 -28 3494
rect -818 3426 -784 3429
rect -62 3426 -28 3450
rect -818 3395 -784 3426
rect -62 3416 -48 3426
rect -48 3416 -28 3426
rect -62 3358 -28 3378
rect -818 3324 -784 3357
rect -62 3344 -48 3358
rect -48 3344 -28 3358
rect -818 3323 -784 3324
rect -62 3290 -28 3306
rect -818 3256 -784 3285
rect -62 3272 -48 3290
rect -48 3272 -28 3290
rect -818 3251 -784 3256
rect -62 3222 -28 3234
rect -818 3188 -784 3213
rect -62 3200 -48 3222
rect -48 3200 -28 3222
rect -818 3179 -784 3188
rect -818 3120 -784 3141
rect -44 3120 -14 3151
rect -14 3120 -10 3151
rect -818 3107 -784 3120
rect -44 3117 -10 3120
rect -818 3052 -784 3069
rect -44 3052 -14 3079
rect -14 3052 -10 3079
rect -818 3035 -784 3052
rect -44 3045 -10 3052
rect -818 2984 -784 2997
rect -44 2984 -14 3007
rect -14 2984 -10 3007
rect -818 2963 -784 2984
rect -44 2973 -10 2984
rect -818 2916 -784 2925
rect -44 2916 -14 2935
rect -14 2916 -10 2935
rect -818 2891 -784 2916
rect -44 2901 -10 2916
rect -818 2848 -784 2853
rect -44 2848 -14 2863
rect -14 2848 -10 2863
rect -818 2819 -784 2848
rect -44 2829 -10 2848
rect -818 2780 -784 2781
rect -44 2780 -14 2791
rect -14 2780 -10 2791
rect -818 2747 -784 2780
rect -44 2757 -10 2780
rect -44 2712 -14 2719
rect -14 2712 -10 2719
rect -818 2678 -784 2709
rect -44 2685 -10 2712
rect -818 2675 -784 2678
rect -44 2644 -14 2647
rect -14 2644 -10 2647
rect -818 2610 -784 2637
rect -44 2613 -10 2644
rect -818 2603 -784 2610
rect -818 2542 -784 2565
rect -44 2542 -10 2575
rect -818 2531 -784 2542
rect -44 2541 -14 2542
rect -14 2541 -10 2542
rect -818 2473 -784 2493
rect -44 2473 -10 2503
rect -818 2459 -784 2473
rect -44 2469 -14 2473
rect -14 2469 -10 2473
rect -818 2404 -784 2421
rect -44 2404 -10 2431
rect -818 2387 -784 2404
rect -44 2397 -14 2404
rect -14 2397 -10 2404
rect -818 2335 -784 2349
rect -44 2335 -10 2359
rect -818 2315 -784 2335
rect -44 2325 -14 2335
rect -14 2325 -10 2335
rect -818 2266 -784 2277
rect -44 2266 -10 2287
rect -818 2243 -784 2266
rect -44 2253 -14 2266
rect -14 2253 -10 2266
rect -818 2197 -784 2205
rect -44 2197 -10 2215
rect -818 2171 -784 2197
rect -44 2181 -14 2197
rect -14 2181 -10 2197
rect -818 2128 -784 2133
rect -44 2128 -10 2143
rect -818 2099 -784 2128
rect -44 2109 -14 2128
rect -14 2109 -10 2128
rect -818 2059 -784 2061
rect -44 2059 -10 2071
rect -818 2027 -784 2059
rect -44 2037 -14 2059
rect -14 2037 -10 2059
rect -44 1990 -10 1999
rect -818 1956 -784 1989
rect -44 1965 -14 1990
rect -14 1965 -10 1990
rect -818 1955 -784 1956
rect -44 1921 -10 1927
rect -818 1887 -784 1917
rect -44 1893 -14 1921
rect -14 1893 -10 1921
rect -818 1883 -784 1887
rect -44 1852 -10 1855
rect -818 1818 -784 1845
rect -44 1821 -14 1852
rect -14 1821 -10 1852
rect -818 1811 -784 1818
rect -818 1749 -784 1773
rect -44 1749 -14 1783
rect -14 1749 -10 1783
rect -818 1739 -784 1749
rect -818 1680 -784 1701
rect -44 1680 -14 1711
rect -14 1680 -10 1711
rect -818 1667 -784 1680
rect -44 1677 -10 1680
rect -818 1611 -784 1629
rect -44 1611 -14 1639
rect -14 1611 -10 1639
rect -818 1595 -784 1611
rect -44 1605 -10 1611
rect -818 1542 -784 1557
rect -44 1542 -14 1567
rect -14 1542 -10 1567
rect -818 1523 -784 1542
rect -44 1533 -10 1542
rect -818 1473 -784 1485
rect -44 1473 -14 1495
rect -14 1473 -10 1495
rect -818 1451 -784 1473
rect -44 1461 -10 1473
rect -818 1404 -784 1413
rect -44 1404 -14 1423
rect -14 1404 -10 1423
rect -818 1379 -784 1404
rect -44 1389 -10 1404
rect -818 1335 -784 1341
rect -44 1335 -14 1351
rect -14 1335 -10 1351
rect -818 1307 -784 1335
rect -44 1317 -10 1335
rect -818 1266 -784 1269
rect -44 1266 -14 1279
rect -14 1266 -10 1279
rect -818 1235 -784 1266
rect -44 1245 -10 1266
rect -44 1197 -14 1207
rect -14 1197 -10 1207
rect -818 1163 -784 1197
rect -44 1173 -10 1197
rect -44 1128 -14 1135
rect -14 1128 -10 1135
rect -818 1093 -784 1125
rect -44 1101 -10 1128
rect -818 1091 -784 1093
rect -44 1059 -14 1063
rect -14 1059 -10 1063
rect -818 1024 -784 1053
rect -44 1029 -10 1059
rect -818 1019 -784 1024
rect -818 955 -784 981
rect -44 956 -10 990
rect -818 947 -784 955
rect -818 886 -784 909
rect -44 886 -10 917
rect -818 875 -784 886
rect -44 883 -14 886
rect -14 883 -10 886
rect -818 817 -784 837
rect -44 817 -10 844
rect -818 803 -784 817
rect -44 810 -14 817
rect -14 810 -10 817
rect -818 748 -784 765
rect -44 748 -10 771
rect -818 731 -784 748
rect -44 737 -14 748
rect -14 737 -10 748
rect -818 679 -784 693
rect -44 679 -10 698
rect -818 659 -784 679
rect -44 664 -14 679
rect -14 664 -10 679
rect -818 610 -784 621
rect -44 610 -10 625
rect -818 587 -784 610
rect -44 591 -14 610
rect -14 591 -10 610
rect -818 541 -784 548
rect -44 541 -10 552
rect -818 514 -784 541
rect -44 518 -14 541
rect -14 518 -10 541
rect -818 472 -784 475
rect -44 472 -10 479
rect -818 441 -784 472
rect -44 445 -14 472
rect -14 445 -10 472
rect -44 403 -10 406
rect -818 369 -784 402
rect -44 372 -14 403
rect -14 372 -10 403
rect -818 368 -784 369
rect -818 300 -784 329
rect -44 300 -14 333
rect -14 300 -10 333
rect -818 295 -784 300
rect -44 299 -10 300
rect -818 231 -784 256
rect -44 231 -14 260
rect -14 231 -10 260
rect -818 222 -784 231
rect -44 226 -10 231
rect -818 162 -784 183
rect -44 162 -14 187
rect -14 162 -10 187
rect -818 149 -784 162
rect -44 153 -10 162
rect 231 4808 265 4842
rect 303 4822 337 4842
rect 303 4808 312 4822
rect 312 4808 337 4822
rect 375 4822 409 4842
rect 375 4808 391 4822
rect 391 4808 409 4822
rect 447 4808 481 4842
rect 519 4822 553 4842
rect 519 4808 525 4822
rect 525 4808 553 4822
rect 171 4744 205 4778
rect 651 4764 662 4782
rect 662 4764 685 4782
rect 171 4668 205 4702
rect 651 4748 685 4764
rect 171 4592 205 4626
rect 284 4625 288 4658
rect 288 4625 318 4658
rect 284 4624 318 4625
rect 284 4556 288 4583
rect 288 4556 318 4583
rect 171 4516 205 4550
rect 284 4549 318 4556
rect 284 4487 288 4508
rect 288 4487 318 4508
rect 284 4474 318 4487
rect 171 4440 205 4474
rect 284 4418 288 4433
rect 288 4418 318 4433
rect 284 4399 318 4418
rect 171 4364 205 4398
rect 284 4349 288 4357
rect 288 4349 318 4357
rect 284 4323 318 4349
rect 171 4288 205 4322
rect 284 4280 288 4281
rect 288 4280 318 4281
rect 284 4247 318 4280
rect 171 4212 205 4246
rect 284 4176 318 4205
rect 284 4171 288 4176
rect 288 4171 318 4176
rect 171 4136 205 4170
rect 284 4107 318 4129
rect 284 4095 288 4107
rect 288 4095 318 4107
rect 171 4059 205 4093
rect 284 4038 318 4053
rect 284 4019 288 4038
rect 288 4019 318 4038
rect 171 3982 205 4016
rect 284 3969 318 3977
rect 284 3943 288 3969
rect 288 3943 318 3969
rect 171 3905 205 3939
rect 284 3900 318 3901
rect 284 3867 288 3900
rect 288 3867 318 3900
rect 171 3828 205 3862
rect 284 3797 288 3825
rect 288 3797 318 3825
rect 284 3791 318 3797
rect 171 3751 205 3785
rect 171 3674 205 3708
rect 171 3597 205 3631
rect 167 3515 201 3549
rect 255 3521 288 3549
rect 288 3521 289 3549
rect 255 3515 289 3521
rect 167 3442 201 3476
rect 255 3452 288 3475
rect 288 3452 289 3475
rect 255 3441 289 3452
rect 167 3370 201 3404
rect 255 3383 288 3401
rect 288 3383 289 3401
rect 255 3367 289 3383
rect 167 3298 201 3332
rect 255 3314 288 3327
rect 288 3314 289 3327
rect 255 3293 289 3314
rect 167 3226 201 3260
rect 255 3245 288 3253
rect 288 3245 289 3253
rect 255 3219 289 3245
rect 167 3154 201 3188
rect 255 3176 288 3179
rect 288 3176 289 3179
rect 255 3145 289 3176
rect 167 3082 201 3116
rect 255 3072 289 3105
rect 255 3071 288 3072
rect 288 3071 289 3072
rect 167 3010 201 3044
rect 255 3003 289 3031
rect 255 2997 288 3003
rect 288 2997 289 3003
rect 167 2938 201 2972
rect 255 2934 289 2957
rect 255 2923 288 2934
rect 288 2923 289 2934
rect 167 2866 201 2900
rect 255 2865 289 2883
rect 255 2849 288 2865
rect 288 2849 289 2865
rect 167 2794 201 2828
rect 255 2796 289 2809
rect 255 2775 288 2796
rect 288 2775 289 2796
rect 167 2722 201 2756
rect 255 2727 289 2735
rect 255 2701 288 2727
rect 288 2701 289 2727
rect 167 2650 201 2684
rect 255 2658 289 2661
rect 255 2627 288 2658
rect 288 2627 289 2658
rect 167 2578 201 2612
rect 255 2555 288 2587
rect 288 2555 289 2587
rect 255 2553 289 2555
rect 167 2506 201 2540
rect 255 2486 288 2514
rect 288 2486 289 2514
rect 255 2480 289 2486
rect 167 2434 201 2468
rect 255 2417 288 2441
rect 288 2417 289 2441
rect 255 2407 289 2417
rect 167 2362 201 2396
rect 255 2348 288 2368
rect 288 2348 289 2368
rect 255 2334 289 2348
rect 167 2290 201 2324
rect 255 2279 288 2295
rect 288 2279 289 2295
rect 255 2261 289 2279
rect 167 2218 201 2252
rect 255 2210 288 2222
rect 288 2210 289 2222
rect 255 2188 289 2210
rect 167 2146 201 2180
rect 255 2141 288 2149
rect 288 2141 289 2149
rect 255 2115 289 2141
rect 167 2074 201 2108
rect 255 2072 288 2076
rect 288 2072 289 2076
rect 255 2042 289 2072
rect 167 2002 201 2036
rect 255 1969 289 2003
rect 167 1930 201 1964
rect 255 1899 289 1930
rect 255 1896 288 1899
rect 288 1896 289 1899
rect 167 1858 201 1892
rect 255 1830 289 1857
rect 255 1823 288 1830
rect 288 1823 289 1830
rect 167 1786 201 1820
rect 255 1761 289 1784
rect 255 1750 288 1761
rect 288 1750 289 1761
rect 167 1714 201 1748
rect 255 1692 289 1711
rect 255 1677 288 1692
rect 288 1677 289 1692
rect 167 1642 201 1676
rect 255 1623 289 1638
rect 255 1604 288 1623
rect 288 1604 289 1623
rect 167 1570 201 1604
rect 255 1554 289 1565
rect 167 1498 201 1532
rect 255 1531 288 1554
rect 288 1531 289 1554
rect 255 1485 289 1492
rect 167 1426 201 1460
rect 255 1458 288 1485
rect 288 1458 289 1485
rect 255 1416 289 1419
rect 167 1354 201 1388
rect 255 1385 288 1416
rect 288 1385 289 1416
rect 167 1282 201 1316
rect 255 1313 288 1346
rect 288 1313 289 1346
rect 255 1312 289 1313
rect 255 1244 288 1273
rect 288 1244 289 1273
rect 167 1210 201 1244
rect 255 1239 289 1244
rect 255 1175 288 1200
rect 288 1175 289 1200
rect 167 1138 201 1172
rect 255 1166 289 1175
rect 255 1106 288 1127
rect 288 1106 289 1127
rect 167 1066 201 1100
rect 255 1093 289 1106
rect 255 1037 288 1054
rect 288 1037 289 1054
rect 167 994 201 1028
rect 255 1020 289 1037
rect 255 968 288 981
rect 288 968 289 981
rect 167 922 201 956
rect 255 947 289 968
rect 255 899 288 908
rect 288 899 289 908
rect 167 850 201 884
rect 255 874 289 899
rect 255 830 288 835
rect 288 830 289 835
rect 167 778 201 812
rect 255 801 289 830
rect 255 761 288 762
rect 288 761 289 762
rect 167 706 201 740
rect 255 728 289 761
rect 167 634 201 668
rect 255 657 289 689
rect 255 655 288 657
rect 288 655 289 657
rect 167 562 201 596
rect 255 588 289 616
rect 255 582 288 588
rect 288 582 289 588
rect 167 490 201 524
rect 255 519 289 543
rect 255 509 288 519
rect 288 509 289 519
rect 167 418 201 452
rect 255 450 289 470
rect 255 436 288 450
rect 288 436 289 450
rect 255 381 289 397
rect 167 346 201 380
rect 255 363 288 381
rect 288 363 289 381
rect 651 4695 662 4708
rect 662 4695 685 4708
rect 651 4674 685 4695
rect 539 4634 573 4658
rect 539 4624 546 4634
rect 546 4624 573 4634
rect 651 4626 662 4634
rect 662 4626 685 4634
rect 651 4600 685 4626
rect 539 4566 573 4583
rect 539 4549 546 4566
rect 546 4549 573 4566
rect 651 4557 662 4561
rect 662 4557 685 4561
rect 651 4527 685 4557
rect 539 4498 573 4508
rect 539 4474 546 4498
rect 546 4474 573 4498
rect 651 4454 685 4488
rect 539 4430 573 4433
rect 539 4399 546 4430
rect 546 4399 573 4430
rect 651 4384 685 4415
rect 651 4381 662 4384
rect 662 4381 685 4384
rect 539 4328 546 4357
rect 546 4328 573 4357
rect 539 4323 573 4328
rect 651 4315 685 4342
rect 651 4308 662 4315
rect 662 4308 685 4315
rect 539 4260 546 4281
rect 546 4260 573 4281
rect 539 4247 573 4260
rect 651 4246 685 4269
rect 651 4235 662 4246
rect 662 4235 685 4246
rect 539 4192 546 4205
rect 546 4192 573 4205
rect 539 4171 573 4192
rect 651 4177 685 4196
rect 651 4162 662 4177
rect 662 4162 685 4177
rect 539 4124 546 4129
rect 546 4124 573 4129
rect 539 4095 573 4124
rect 651 4108 685 4123
rect 651 4089 662 4108
rect 662 4089 685 4108
rect 539 4022 573 4053
rect 651 4039 685 4050
rect 539 4019 546 4022
rect 546 4019 573 4022
rect 651 4016 662 4039
rect 662 4016 685 4039
rect 539 3954 573 3977
rect 651 3970 685 3977
rect 539 3943 546 3954
rect 546 3943 573 3954
rect 651 3943 662 3970
rect 662 3943 685 3970
rect 651 3901 685 3904
rect 539 3886 573 3901
rect 539 3867 546 3886
rect 546 3867 573 3886
rect 651 3870 662 3901
rect 662 3870 685 3901
rect 539 3818 573 3825
rect 539 3791 546 3818
rect 546 3791 573 3818
rect 651 3798 662 3831
rect 662 3798 685 3831
rect 651 3797 685 3798
rect 651 3729 662 3758
rect 662 3729 685 3758
rect 370 3660 404 3694
rect 651 3724 685 3729
rect 370 3587 404 3621
rect 370 3547 404 3548
rect 370 3514 404 3547
rect 370 3445 404 3475
rect 370 3441 404 3445
rect 370 3377 404 3402
rect 370 3368 404 3377
rect 370 3309 404 3329
rect 370 3295 404 3309
rect 370 3241 404 3256
rect 370 3222 404 3241
rect 370 3173 404 3183
rect 370 3149 404 3173
rect 370 3105 404 3110
rect 370 3076 404 3105
rect 370 3003 404 3037
rect 370 2935 404 2964
rect 370 2930 404 2935
rect 370 2867 404 2891
rect 370 2857 404 2867
rect 370 2799 404 2818
rect 370 2784 404 2799
rect 370 2731 404 2745
rect 370 2711 404 2731
rect 370 2663 404 2673
rect 370 2639 404 2663
rect 370 2567 404 2601
rect 370 2495 404 2529
rect 370 2426 404 2457
rect 370 2423 404 2426
rect 370 2358 404 2385
rect 370 2351 404 2358
rect 370 2290 404 2313
rect 370 2279 404 2290
rect 370 2222 404 2241
rect 370 2207 404 2222
rect 370 2154 404 2169
rect 370 2135 404 2154
rect 370 2086 404 2097
rect 370 2063 404 2086
rect 370 1984 404 2016
rect 370 1982 404 1984
rect 370 1916 404 1943
rect 370 1909 404 1916
rect 370 1848 404 1870
rect 370 1836 404 1848
rect 370 1780 404 1797
rect 370 1763 404 1780
rect 370 1712 404 1725
rect 370 1691 404 1712
rect 370 1644 404 1653
rect 370 1619 404 1644
rect 370 1576 404 1581
rect 370 1547 404 1576
rect 370 1475 404 1509
rect 370 1403 404 1437
rect 472 3640 506 3659
rect 472 3625 506 3640
rect 472 3552 506 3586
rect 472 3479 506 3513
rect 472 3406 506 3440
rect 472 3333 506 3367
rect 472 3260 506 3294
rect 472 3187 506 3221
rect 472 3114 506 3148
rect 472 3040 506 3074
rect 472 2966 506 3000
rect 472 2892 506 2926
rect 472 2818 506 2852
rect 472 2744 506 2778
rect 472 2670 506 2704
rect 472 2596 506 2630
rect 472 2553 506 2556
rect 472 2522 506 2553
rect 472 2448 506 2482
rect 472 2374 506 2408
rect 472 2300 506 2334
rect 472 2226 506 2260
rect 472 2152 506 2186
rect 472 2078 506 2112
rect 472 2004 506 2038
rect 472 1930 506 1964
rect 472 1856 506 1890
rect 472 1782 506 1816
rect 472 1708 506 1742
rect 472 1634 506 1668
rect 472 1560 506 1594
rect 472 1486 506 1520
rect 472 1434 506 1446
rect 472 1412 506 1434
rect 651 3660 662 3685
rect 662 3660 685 3685
rect 651 3651 685 3660
rect 651 3591 662 3612
rect 662 3591 685 3612
rect 651 3578 685 3591
rect 651 3522 662 3539
rect 662 3522 685 3539
rect 651 3505 685 3522
rect 651 3453 662 3466
rect 662 3453 685 3466
rect 651 3432 685 3453
rect 651 3384 662 3393
rect 662 3384 685 3393
rect 651 3359 685 3384
rect 651 3315 662 3320
rect 662 3315 685 3320
rect 651 3286 685 3315
rect 651 3246 662 3247
rect 662 3246 685 3247
rect 651 3213 685 3246
rect 651 3142 685 3174
rect 651 3140 662 3142
rect 662 3140 685 3142
rect 651 3073 685 3101
rect 651 3067 662 3073
rect 662 3067 685 3073
rect 651 3004 685 3028
rect 651 2994 662 3004
rect 662 2994 685 3004
rect 651 2935 685 2955
rect 651 2921 662 2935
rect 662 2921 685 2935
rect 651 2866 685 2882
rect 651 2848 662 2866
rect 662 2848 685 2866
rect 651 2797 685 2809
rect 651 2775 662 2797
rect 662 2775 685 2797
rect 651 2728 685 2736
rect 651 2702 662 2728
rect 662 2702 685 2728
rect 651 2659 685 2663
rect 651 2629 662 2659
rect 662 2629 685 2659
rect 651 2556 662 2590
rect 662 2556 685 2590
rect 651 2487 662 2517
rect 662 2487 685 2517
rect 651 2483 685 2487
rect 651 2418 662 2444
rect 662 2418 685 2444
rect 651 2410 685 2418
rect 651 2349 662 2371
rect 662 2349 685 2371
rect 651 2337 685 2349
rect 651 2280 662 2298
rect 662 2280 685 2298
rect 651 2264 685 2280
rect 651 2211 662 2225
rect 662 2211 685 2225
rect 651 2191 685 2211
rect 651 2142 662 2152
rect 662 2142 685 2152
rect 651 2118 685 2142
rect 651 2073 662 2079
rect 662 2073 685 2079
rect 651 2045 685 2073
rect 668 1900 702 1924
rect 668 1890 696 1900
rect 696 1890 702 1900
rect 756 1890 790 1924
rect 668 1831 702 1852
rect 668 1818 696 1831
rect 696 1818 702 1831
rect 756 1817 790 1851
rect 668 1762 702 1780
rect 668 1746 696 1762
rect 696 1746 702 1762
rect 756 1744 790 1778
rect 668 1693 702 1708
rect 668 1674 696 1693
rect 696 1674 702 1693
rect 756 1671 790 1705
rect 668 1624 702 1636
rect 668 1602 696 1624
rect 696 1602 702 1624
rect 756 1598 790 1632
rect 668 1555 702 1564
rect 668 1530 696 1555
rect 696 1530 702 1555
rect 756 1525 790 1559
rect 668 1486 702 1492
rect 668 1458 696 1486
rect 696 1458 702 1486
rect 756 1452 790 1486
rect 668 1417 702 1419
rect 370 1331 404 1365
rect 668 1385 696 1417
rect 696 1385 702 1417
rect 756 1379 790 1413
rect 370 1292 404 1293
rect 370 1259 404 1292
rect 370 1190 404 1221
rect 370 1187 404 1190
rect 370 1122 404 1149
rect 370 1115 404 1122
rect 370 1054 404 1077
rect 370 1043 404 1054
rect 370 986 404 1005
rect 370 971 404 986
rect 370 918 404 933
rect 370 899 404 918
rect 370 850 404 861
rect 370 827 404 850
rect 370 782 404 789
rect 370 755 404 782
rect 370 714 404 717
rect 370 683 404 714
rect 370 612 404 645
rect 370 611 404 612
rect 370 544 404 573
rect 370 539 404 544
rect 370 476 404 501
rect 370 467 404 476
rect 668 1314 696 1346
rect 696 1314 702 1346
rect 668 1312 702 1314
rect 756 1306 790 1340
rect 668 1245 696 1273
rect 696 1245 702 1273
rect 668 1239 702 1245
rect 756 1233 790 1267
rect 668 1176 696 1200
rect 696 1176 702 1200
rect 668 1166 702 1176
rect 756 1160 790 1194
rect 668 1107 696 1127
rect 696 1107 702 1127
rect 668 1093 702 1107
rect 756 1087 790 1121
rect 668 1038 696 1054
rect 696 1038 702 1054
rect 668 1020 702 1038
rect 756 1014 790 1048
rect 668 969 696 981
rect 696 969 702 981
rect 668 947 702 969
rect 756 940 790 974
rect 668 900 696 908
rect 696 900 702 908
rect 668 874 702 900
rect 756 866 790 900
rect 668 831 696 835
rect 696 831 702 835
rect 668 801 702 831
rect 756 792 790 826
rect 668 728 702 762
rect 756 718 790 752
rect 668 658 702 689
rect 668 655 696 658
rect 696 655 702 658
rect 756 644 790 678
rect 668 589 702 616
rect 668 582 696 589
rect 696 582 702 589
rect 756 570 790 604
rect 668 520 702 543
rect 668 509 696 520
rect 696 509 702 520
rect 756 496 790 530
rect 668 451 702 470
rect 668 436 696 451
rect 696 436 702 451
rect 756 422 790 456
rect 668 382 702 397
rect 668 363 696 382
rect 696 363 702 382
rect 756 348 790 382
rect 255 312 289 324
rect 167 274 201 308
rect 255 290 288 312
rect 288 290 289 312
rect 338 290 372 324
rect 421 290 455 324
rect 504 290 538 324
rect 586 290 620 324
rect 668 290 702 324
rect 756 274 790 308
rect 239 202 273 236
rect 313 202 347 236
rect 387 202 421 236
rect 461 202 495 236
rect 535 202 569 236
rect 609 202 643 236
rect 683 202 717 236
rect -818 93 -784 110
rect -44 93 -14 114
rect -14 93 -10 114
rect -818 76 -784 93
rect -44 80 -10 93
rect 59 68 92 95
rect 92 68 93 95
rect 134 68 161 95
rect 161 68 168 95
rect 209 68 230 95
rect 230 68 243 95
rect 284 68 300 95
rect 300 68 318 95
rect 359 68 370 95
rect 370 68 393 95
rect 434 68 440 95
rect 440 68 468 95
rect 509 68 510 95
rect 510 68 543 95
rect 584 68 614 95
rect 614 68 618 95
rect 659 68 684 95
rect 684 68 693 95
rect 734 68 754 95
rect 754 68 768 95
rect 808 68 824 95
rect 824 68 842 95
rect 59 61 93 68
rect 134 61 168 68
rect 209 61 243 68
rect 284 61 318 68
rect 359 61 393 68
rect 434 61 468 68
rect 509 61 543 68
rect 584 61 618 68
rect 659 61 693 68
rect 734 61 768 68
rect 808 61 842 68
rect -818 24 -784 37
rect -44 24 -14 41
rect -14 24 -10 41
rect -818 3 -784 24
rect -44 7 -10 24
rect 36 -15 70 19
rect 113 0 126 19
rect 126 0 147 19
rect 190 0 195 19
rect 195 0 224 19
rect 267 0 300 19
rect 300 0 301 19
rect 344 0 370 19
rect 370 0 378 19
rect 421 0 440 19
rect 440 0 455 19
rect 498 0 510 19
rect 510 0 532 19
rect 575 0 580 19
rect 580 0 609 19
rect 653 0 684 19
rect 684 0 687 19
rect 731 0 754 19
rect 754 0 765 19
rect 809 0 824 19
rect 824 0 843 19
rect 113 -15 147 0
rect 190 -15 224 0
rect 267 -15 301 0
rect 344 -15 378 0
rect 421 -15 455 0
rect 498 -15 532 0
rect 575 -15 609 0
rect 653 -15 687 0
rect 731 -15 765 0
rect 809 -15 843 0
rect -818 -68 -784 -36
rect -818 -70 -784 -68
rect 36 -99 70 -65
rect 113 -68 140 -65
rect 140 -68 147 -65
rect 190 -68 209 -65
rect 209 -68 224 -65
rect 267 -68 278 -65
rect 278 -68 301 -65
rect 344 -68 347 -65
rect 347 -68 378 -65
rect 421 -68 450 -65
rect 450 -68 455 -65
rect 498 -68 519 -65
rect 519 -68 532 -65
rect 575 -68 588 -65
rect 588 -68 609 -65
rect 653 -68 657 -65
rect 657 -68 687 -65
rect 731 -68 761 -65
rect 761 -68 765 -65
rect 809 -68 830 -65
rect 830 -68 843 -65
rect 113 -99 147 -68
rect 190 -99 224 -68
rect 267 -99 301 -68
rect 344 -99 378 -68
rect 421 -99 455 -68
rect 498 -99 532 -68
rect 575 -99 609 -68
rect 653 -99 687 -68
rect 731 -99 765 -68
rect 809 -99 843 -68
rect -818 -139 -784 -109
rect -818 -143 -784 -139
rect -818 -210 -784 -182
rect 36 -183 70 -149
rect 113 -176 147 -149
rect 190 -176 224 -149
rect 267 -176 301 -149
rect 344 -176 378 -149
rect 421 -176 455 -149
rect 498 -176 532 -149
rect 575 -176 609 -149
rect 653 -176 687 -149
rect 731 -176 765 -149
rect 809 -176 843 -149
rect 113 -183 140 -176
rect 140 -183 147 -176
rect 190 -183 209 -176
rect 209 -183 224 -176
rect 267 -183 278 -176
rect 278 -183 301 -176
rect 344 -183 347 -176
rect 347 -183 378 -176
rect 421 -183 450 -176
rect 450 -183 455 -176
rect 498 -183 519 -176
rect 519 -183 532 -176
rect 575 -183 588 -176
rect 588 -183 609 -176
rect 653 -183 657 -176
rect 657 -183 687 -176
rect 731 -183 761 -176
rect 761 -183 765 -176
rect 809 -183 830 -176
rect 830 -183 843 -176
rect -818 -216 -784 -210
rect -42 -247 -8 -215
rect -818 -281 -784 -255
rect -730 -281 -716 -255
rect -716 -281 -696 -255
rect -42 -249 -33 -247
rect -33 -249 -8 -247
rect 36 -267 70 -233
rect 113 -247 147 -233
rect 190 -247 224 -233
rect 267 -247 301 -233
rect 344 -247 378 -233
rect 421 -247 455 -233
rect 498 -247 532 -233
rect 575 -247 609 -233
rect 653 -247 687 -233
rect 731 -247 765 -233
rect 809 -247 843 -233
rect 113 -267 140 -247
rect 140 -267 147 -247
rect 190 -267 209 -247
rect 209 -267 224 -247
rect 267 -267 278 -247
rect 278 -267 301 -247
rect 344 -267 347 -247
rect 347 -267 378 -247
rect 421 -267 450 -247
rect 450 -267 455 -247
rect 498 -267 519 -247
rect 519 -267 532 -247
rect 575 -267 588 -247
rect 588 -267 609 -247
rect 653 -267 657 -247
rect 657 -267 687 -247
rect 731 -267 761 -247
rect 761 -267 765 -247
rect 809 -267 830 -247
rect 830 -267 843 -247
rect -818 -289 -784 -281
rect -730 -289 -696 -281
rect -114 -318 -80 -287
rect -42 -318 -8 -287
rect -730 -352 -716 -327
rect -716 -352 -696 -327
rect -114 -321 -102 -318
rect -102 -321 -80 -318
rect -42 -321 -33 -318
rect -33 -321 -8 -318
rect 36 -351 70 -317
rect 113 -318 147 -317
rect 190 -318 224 -317
rect 267 -318 301 -317
rect 344 -318 378 -317
rect 421 -318 455 -317
rect 498 -318 532 -317
rect 575 -318 609 -317
rect 653 -318 687 -317
rect 731 -318 765 -317
rect 809 -318 843 -317
rect 113 -351 140 -318
rect 140 -351 147 -318
rect 190 -351 209 -318
rect 209 -351 224 -318
rect 267 -351 278 -318
rect 278 -351 301 -318
rect 344 -351 347 -318
rect 347 -351 378 -318
rect 421 -351 450 -318
rect 450 -351 455 -318
rect 498 -351 519 -318
rect 519 -351 532 -318
rect 575 -351 588 -318
rect 588 -351 609 -318
rect 653 -351 657 -318
rect 657 -351 687 -318
rect 731 -351 761 -318
rect 761 -351 765 -318
rect 809 -351 830 -318
rect 830 -351 843 -318
rect -730 -361 -696 -352
<< metal1 >>
rect -824 14517 -778 14529
rect -824 14483 -818 14517
rect -784 14483 -778 14517
rect -824 14445 -778 14483
rect -824 14411 -818 14445
rect -784 14411 -778 14445
rect -824 14373 -778 14411
rect -824 14339 -818 14373
rect -784 14339 -778 14373
rect -824 14301 -778 14339
rect -824 14267 -818 14301
rect -784 14267 -778 14301
rect -824 14229 -778 14267
rect -824 14195 -818 14229
rect -784 14195 -778 14229
rect -824 14157 -778 14195
rect -824 14123 -818 14157
rect -784 14123 -778 14157
rect -824 14085 -778 14123
rect -824 14051 -818 14085
rect -784 14051 -778 14085
tri -826 14039 -824 14041 se
rect -824 14039 -778 14051
tri -830 14035 -826 14039 se
rect -826 14035 -778 14039
rect -830 14029 -778 14035
rect -830 13955 -778 13977
rect -830 13881 -778 13903
rect -830 13807 -778 13829
rect -830 13733 -778 13755
rect -830 13675 -778 13681
tri -830 13669 -824 13675 ne
rect -824 13653 -778 13675
rect -824 13619 -818 13653
rect -784 13619 -778 13653
rect -824 13581 -778 13619
rect -824 13547 -818 13581
rect -784 13547 -778 13581
rect -824 13509 -778 13547
rect -824 13475 -818 13509
rect -784 13475 -778 13509
rect -824 13437 -778 13475
rect -824 13403 -818 13437
rect -784 13403 -778 13437
rect -824 13365 -778 13403
rect -824 13331 -818 13365
rect -784 13331 -778 13365
rect -824 13293 -778 13331
rect -824 13259 -818 13293
rect -784 13259 -778 13293
rect -824 13221 -778 13259
rect -824 13187 -818 13221
rect -784 13187 -778 13221
rect -824 13149 -778 13187
rect -824 13115 -818 13149
rect -784 13115 -778 13149
rect -824 13077 -778 13115
rect -824 13043 -818 13077
rect -784 13043 -778 13077
rect -824 13005 -778 13043
rect -824 12971 -818 13005
rect -784 12971 -778 13005
rect -824 12933 -778 12971
rect -824 12899 -818 12933
rect -784 12899 -778 12933
rect -824 12861 -778 12899
rect -824 12827 -818 12861
rect -784 12827 -778 12861
rect -824 12789 -778 12827
rect -824 12755 -818 12789
rect -784 12755 -778 12789
rect -824 12717 -778 12755
rect -824 12683 -818 12717
rect -784 12683 -778 12717
rect -824 12645 -778 12683
rect -824 12611 -818 12645
rect -784 12611 -778 12645
rect -824 12573 -778 12611
rect -824 12539 -818 12573
rect -784 12539 -778 12573
rect -824 12501 -778 12539
rect -824 12467 -818 12501
rect -784 12467 -778 12501
rect -824 12429 -778 12467
rect -824 12395 -818 12429
rect -784 12395 -778 12429
rect -824 12357 -778 12395
rect -824 12323 -818 12357
rect -784 12323 -778 12357
rect -824 12285 -778 12323
rect -824 12251 -818 12285
rect -784 12251 -778 12285
rect -824 12213 -778 12251
rect -824 12179 -818 12213
rect -784 12179 -778 12213
rect -824 12141 -778 12179
rect -824 12107 -818 12141
rect -784 12107 -778 12141
rect -824 12069 -778 12107
rect -824 12035 -818 12069
rect -784 12035 -778 12069
rect -824 11997 -778 12035
rect -824 11963 -818 11997
rect -784 11963 -778 11997
rect -824 11925 -778 11963
rect -824 11891 -818 11925
rect -784 11891 -778 11925
rect -824 11853 -778 11891
rect -824 11819 -818 11853
rect -784 11819 -778 11853
rect -824 11781 -778 11819
rect -824 11747 -818 11781
rect -784 11747 -778 11781
rect -824 11709 -778 11747
rect -824 11675 -818 11709
rect -784 11675 -778 11709
rect -824 11637 -778 11675
rect -824 11603 -818 11637
rect -784 11603 -778 11637
rect -824 11565 -778 11603
rect -824 11531 -818 11565
rect -784 11531 -778 11565
rect -824 11493 -778 11531
rect -824 11459 -818 11493
rect -784 11459 -778 11493
rect -824 11421 -778 11459
rect -824 11387 -818 11421
rect -784 11387 -778 11421
rect -824 11349 -778 11387
rect -824 11315 -818 11349
rect -784 11315 -778 11349
rect -824 11277 -778 11315
rect -824 11243 -818 11277
rect -784 11243 -778 11277
rect -824 11205 -778 11243
rect -824 11171 -818 11205
rect -784 11171 -778 11205
rect -824 11133 -778 11171
rect -824 11099 -818 11133
rect -784 11099 -778 11133
rect -824 11061 -778 11099
rect -824 11027 -818 11061
rect -784 11027 -778 11061
rect -824 10989 -778 11027
rect -824 10955 -818 10989
rect -784 10955 -778 10989
rect -824 10917 -778 10955
rect -824 10883 -818 10917
rect -784 10883 -778 10917
rect -824 10845 -778 10883
rect -824 10811 -818 10845
rect -784 10811 -778 10845
rect -824 10773 -778 10811
rect -824 10739 -818 10773
rect -784 10739 -778 10773
rect -824 10701 -778 10739
rect -824 10667 -818 10701
rect -784 10667 -778 10701
rect -824 10629 -778 10667
rect -824 10595 -818 10629
rect -784 10595 -778 10629
rect -824 10557 -778 10595
rect -824 10523 -818 10557
rect -784 10523 -778 10557
rect -824 10485 -778 10523
rect -824 10451 -818 10485
rect -784 10451 -778 10485
rect -824 10413 -778 10451
rect -824 10379 -818 10413
rect -784 10379 -778 10413
rect -824 10341 -778 10379
rect -824 10307 -818 10341
rect -784 10307 -778 10341
rect -824 10269 -778 10307
rect -824 10235 -818 10269
rect -784 10235 -778 10269
rect -824 10197 -778 10235
rect -824 10163 -818 10197
rect -784 10163 -778 10197
rect -824 10125 -778 10163
rect -824 10091 -818 10125
rect -784 10091 -778 10125
rect -824 10053 -778 10091
rect -824 10019 -818 10053
rect -784 10019 -778 10053
rect -824 9981 -778 10019
rect -824 9947 -818 9981
rect -784 9947 -778 9981
rect -824 9909 -778 9947
rect -824 9875 -818 9909
rect -784 9875 -778 9909
rect -824 9837 -778 9875
rect -824 9803 -818 9837
rect -784 9803 -778 9837
rect -824 9765 -778 9803
rect -824 9731 -818 9765
rect -784 9731 -778 9765
rect -824 9693 -778 9731
rect -824 9659 -818 9693
rect -784 9659 -778 9693
rect -824 9621 -778 9659
rect -824 9587 -818 9621
rect -784 9587 -778 9621
rect -824 9549 -778 9587
rect -824 9515 -818 9549
rect -784 9515 -778 9549
rect -824 9477 -778 9515
rect -824 9443 -818 9477
rect -784 9443 -778 9477
rect -824 9405 -778 9443
rect -824 9371 -818 9405
rect -784 9371 -778 9405
rect -824 9333 -778 9371
rect -824 9299 -818 9333
rect -784 9299 -778 9333
rect -824 9261 -778 9299
rect -824 9227 -818 9261
rect -784 9227 -778 9261
rect -824 9189 -778 9227
rect -824 9155 -818 9189
rect -784 9155 -778 9189
rect -824 9117 -778 9155
rect -824 9083 -818 9117
rect -784 9083 -778 9117
rect -824 9045 -778 9083
rect -824 9011 -818 9045
rect -784 9011 -778 9045
rect -824 8973 -778 9011
rect -824 8939 -818 8973
rect -784 8939 -778 8973
rect -824 8901 -778 8939
rect -824 8867 -818 8901
rect -784 8867 -778 8901
rect -824 8829 -778 8867
rect -824 8795 -818 8829
rect -784 8795 -778 8829
rect -824 8757 -778 8795
rect -824 8723 -818 8757
rect -784 8723 -778 8757
rect -824 8685 -778 8723
rect -824 8651 -818 8685
rect -784 8651 -778 8685
rect -824 8613 -778 8651
rect -824 8579 -818 8613
rect -784 8579 -778 8613
rect -824 8541 -778 8579
rect -824 8507 -818 8541
rect -784 8507 -778 8541
rect -824 8469 -778 8507
rect -824 8435 -818 8469
rect -784 8435 -778 8469
rect -824 8397 -778 8435
rect -824 8363 -818 8397
rect -784 8363 -778 8397
rect -824 8325 -778 8363
rect -824 8291 -818 8325
rect -784 8291 -778 8325
rect -824 8253 -778 8291
rect -824 8219 -818 8253
rect -784 8219 -778 8253
rect -824 8181 -778 8219
rect -824 8147 -818 8181
rect -784 8147 -778 8181
rect -824 8109 -778 8147
rect -824 8075 -818 8109
rect -784 8075 -778 8109
rect -824 8037 -778 8075
rect -824 8003 -818 8037
rect -784 8003 -778 8037
rect -824 7965 -778 8003
rect -824 7931 -818 7965
rect -784 7931 -778 7965
rect -824 7893 -778 7931
rect -824 7859 -818 7893
rect -784 7859 -778 7893
rect -824 7821 -778 7859
rect -824 7787 -818 7821
rect -784 7787 -778 7821
rect -824 7749 -778 7787
rect -824 7715 -818 7749
rect -784 7715 -778 7749
rect -824 7677 -778 7715
rect -824 7643 -818 7677
rect -784 7643 -778 7677
rect -824 7605 -778 7643
rect -824 7571 -818 7605
rect -784 7571 -778 7605
rect -824 7533 -778 7571
rect -824 7499 -818 7533
rect -784 7499 -778 7533
rect -824 7461 -778 7499
rect -824 7427 -818 7461
rect -784 7427 -778 7461
rect -824 7389 -778 7427
rect -824 7355 -818 7389
rect -784 7355 -778 7389
rect -824 7317 -778 7355
rect -824 7283 -818 7317
rect -784 7283 -778 7317
rect -824 7245 -778 7283
rect -824 7211 -818 7245
rect -784 7211 -778 7245
rect -824 7173 -778 7211
rect -824 7139 -818 7173
rect -784 7139 -778 7173
rect -824 7101 -778 7139
rect -824 7067 -818 7101
rect -784 7067 -778 7101
rect -824 7029 -778 7067
rect -824 6995 -818 7029
rect -784 6995 -778 7029
rect -824 6957 -778 6995
rect -824 6923 -818 6957
rect -784 6923 -778 6957
rect -824 6885 -778 6923
rect -824 6851 -818 6885
rect -784 6851 -778 6885
rect -824 6813 -778 6851
rect -824 6779 -818 6813
rect -784 6779 -778 6813
rect -824 6741 -778 6779
rect -824 6707 -818 6741
rect -784 6707 -778 6741
rect -824 6669 -778 6707
rect -824 6635 -818 6669
rect -784 6635 -778 6669
rect -824 6597 -778 6635
rect -824 6563 -818 6597
rect -784 6563 -778 6597
rect -824 6525 -778 6563
rect -824 6491 -818 6525
rect -784 6491 -778 6525
rect -824 6453 -778 6491
rect -824 6419 -818 6453
rect -784 6419 -778 6453
rect -824 6381 -778 6419
rect -824 6347 -818 6381
rect -784 6347 -778 6381
rect -824 6309 -778 6347
rect -824 6275 -818 6309
rect -784 6275 -778 6309
rect -824 6237 -778 6275
rect -824 6203 -818 6237
rect -784 6203 -778 6237
rect -824 6165 -778 6203
rect -824 6131 -818 6165
rect -784 6131 -778 6165
rect -824 6093 -778 6131
rect -824 6059 -818 6093
rect -784 6059 -778 6093
rect -824 6021 -778 6059
rect -824 5987 -818 6021
rect -784 5987 -778 6021
rect -824 5949 -778 5987
rect -824 5915 -818 5949
rect -784 5915 -778 5949
rect -824 5877 -778 5915
rect -824 5843 -818 5877
rect -784 5843 -778 5877
rect -824 5805 -778 5843
rect -824 5771 -818 5805
rect -784 5771 -778 5805
rect -824 5733 -778 5771
rect -824 5699 -818 5733
rect -784 5699 -778 5733
rect -824 5661 -778 5699
rect -824 5627 -818 5661
rect -784 5627 -778 5661
rect -824 5589 -778 5627
rect -824 5555 -818 5589
rect -784 5555 -778 5589
rect -824 5517 -778 5555
rect -824 5483 -818 5517
rect -784 5483 -778 5517
rect -824 5445 -778 5483
rect -824 5411 -818 5445
rect -784 5411 -778 5445
rect -824 5373 -778 5411
rect -824 5339 -818 5373
rect -784 5339 -778 5373
rect -824 5301 -778 5339
rect -824 5267 -818 5301
rect -784 5267 -778 5301
rect -824 5229 -778 5267
rect -824 5195 -818 5229
rect -784 5195 -778 5229
rect -824 5157 -778 5195
rect -824 5123 -818 5157
rect -784 5123 -778 5157
rect -824 5085 -778 5123
rect -824 5051 -818 5085
rect -784 5051 -778 5085
rect -824 5013 -778 5051
rect -824 4979 -818 5013
rect -784 4979 -778 5013
rect -824 4941 -778 4979
rect -824 4907 -818 4941
rect -784 4907 -778 4941
rect -824 4869 -778 4907
rect -824 4835 -818 4869
rect -784 4835 -778 4869
rect -824 4797 -778 4835
rect -824 4763 -818 4797
rect -784 4763 -778 4797
rect -824 4725 -778 4763
rect -824 4691 -818 4725
rect -784 4691 -778 4725
rect -824 4653 -778 4691
rect -824 4619 -818 4653
rect -784 4619 -778 4653
rect -824 4581 -778 4619
rect -824 4547 -818 4581
rect -784 4547 -778 4581
rect -824 4509 -778 4547
rect -824 4475 -818 4509
rect -784 4475 -778 4509
rect -824 4437 -778 4475
rect -824 4403 -818 4437
rect -784 4403 -778 4437
rect -824 4365 -778 4403
rect -824 4331 -818 4365
rect -784 4331 -778 4365
rect -824 4293 -778 4331
rect -824 4259 -818 4293
rect -784 4259 -778 4293
rect -824 4221 -778 4259
rect -824 4187 -818 4221
rect -784 4187 -778 4221
rect -824 4149 -778 4187
rect -824 4115 -818 4149
rect -784 4115 -778 4149
rect -824 4077 -778 4115
rect -824 4043 -818 4077
rect -784 4043 -778 4077
rect -824 4005 -778 4043
rect -824 3971 -818 4005
rect -784 3971 -778 4005
rect -824 3933 -778 3971
rect -824 3899 -818 3933
rect -784 3899 -778 3933
rect -824 3861 -778 3899
rect -824 3827 -818 3861
rect -784 3827 -778 3861
rect -824 3789 -778 3827
rect -824 3755 -818 3789
rect -784 3755 -778 3789
rect -824 3717 -778 3755
rect -824 3683 -818 3717
rect -784 3683 -778 3717
rect -824 3645 -778 3683
rect -824 3611 -818 3645
rect -784 3611 -778 3645
rect -824 3573 -778 3611
rect -824 3539 -818 3573
rect -784 3539 -778 3573
rect -824 3501 -778 3539
rect -824 3467 -818 3501
rect -784 3467 -778 3501
rect -824 3429 -778 3467
rect -311 14505 -117 14517
rect -311 14471 -305 14505
rect -271 14471 -231 14505
rect -197 14471 -157 14505
rect -123 14471 -117 14505
rect -311 14433 -117 14471
rect -311 14399 -305 14433
rect -271 14399 -231 14433
rect -197 14399 -157 14433
rect -123 14399 -117 14433
rect -311 14361 -117 14399
rect -311 14327 -305 14361
rect -271 14327 -231 14361
rect -197 14327 -157 14361
rect -123 14327 -117 14361
rect -311 14289 -117 14327
rect -311 14255 -305 14289
rect -271 14255 -231 14289
rect -197 14255 -157 14289
rect -123 14255 -117 14289
rect -311 14217 -117 14255
rect -311 14183 -305 14217
rect -271 14183 -231 14217
rect -197 14183 -157 14217
rect -123 14183 -117 14217
rect -311 14145 -117 14183
rect -311 14111 -305 14145
rect -271 14111 -231 14145
rect -197 14111 -157 14145
rect -123 14111 -117 14145
rect -311 14073 -117 14111
rect -311 14039 -305 14073
rect -271 14039 -231 14073
rect -197 14039 -157 14073
rect -123 14039 -117 14073
rect -311 14027 -117 14039
rect -311 13975 -310 14027
rect -258 13975 -242 14027
rect -190 13975 -174 14027
rect -122 13975 -117 14027
rect -311 13967 -305 13975
rect -271 13967 -231 13975
rect -197 13967 -157 13975
rect -123 13967 -117 13975
rect -311 13930 -117 13967
rect -311 13878 -310 13930
rect -258 13878 -242 13930
rect -190 13878 -174 13930
rect -122 13878 -117 13930
rect -311 13857 -117 13878
rect -311 13833 -305 13857
rect -271 13833 -231 13857
rect -197 13833 -157 13857
rect -123 13833 -117 13857
rect -311 13781 -310 13833
rect -258 13781 -242 13833
rect -190 13781 -174 13833
rect -122 13781 -117 13833
rect -311 13751 -305 13781
rect -271 13751 -231 13781
rect -197 13751 -157 13781
rect -123 13751 -117 13781
rect -311 13735 -117 13751
rect -311 13683 -310 13735
rect -258 13683 -242 13735
rect -190 13683 -174 13735
rect -122 13683 -117 13735
rect -311 13679 -305 13683
rect -271 13679 -231 13683
rect -197 13679 -157 13683
rect -123 13679 -117 13683
rect -311 13641 -117 13679
rect -311 13607 -305 13641
rect -271 13607 -231 13641
rect -197 13607 -157 13641
rect -123 13607 -117 13641
rect -311 13569 -117 13607
rect -311 13535 -305 13569
rect -271 13535 -231 13569
rect -197 13535 -157 13569
rect -123 13535 -117 13569
rect -311 13497 -117 13535
rect -311 13463 -305 13497
rect -271 13463 -231 13497
rect -197 13463 -157 13497
rect -123 13463 -117 13497
rect -311 13425 -117 13463
rect -311 13391 -305 13425
rect -271 13391 -231 13425
rect -197 13391 -157 13425
rect -123 13391 -117 13425
rect -311 13353 -117 13391
rect -311 13319 -305 13353
rect -271 13319 -231 13353
rect -197 13319 -157 13353
rect -123 13319 -117 13353
rect -311 13281 -117 13319
rect -311 13247 -305 13281
rect -271 13247 -231 13281
rect -197 13247 -157 13281
rect -123 13247 -117 13281
rect -311 13209 -117 13247
rect -311 13175 -305 13209
rect -271 13175 -231 13209
rect -197 13175 -157 13209
rect -123 13175 -117 13209
rect -311 13137 -117 13175
rect -311 13103 -305 13137
rect -271 13103 -231 13137
rect -197 13103 -157 13137
rect -123 13103 -117 13137
rect -311 13065 -117 13103
rect -311 13031 -305 13065
rect -271 13031 -231 13065
rect -197 13031 -157 13065
rect -123 13031 -117 13065
rect -311 12993 -117 13031
rect -311 12959 -305 12993
rect -271 12959 -231 12993
rect -197 12959 -157 12993
rect -123 12959 -117 12993
rect -311 12921 -117 12959
rect -311 12887 -305 12921
rect -271 12887 -231 12921
rect -197 12887 -157 12921
rect -123 12887 -117 12921
rect -311 12849 -117 12887
rect -311 12815 -305 12849
rect -271 12815 -231 12849
rect -197 12815 -157 12849
rect -123 12815 -117 12849
rect -311 12777 -117 12815
rect -311 12743 -305 12777
rect -271 12743 -231 12777
rect -197 12743 -157 12777
rect -123 12743 -117 12777
rect -311 12705 -117 12743
rect -311 12671 -305 12705
rect -271 12671 -231 12705
rect -197 12671 -157 12705
rect -123 12671 -117 12705
rect -311 12633 -117 12671
rect -311 12599 -305 12633
rect -271 12599 -231 12633
rect -197 12599 -157 12633
rect -123 12599 -117 12633
rect -311 12561 -117 12599
rect -311 12527 -305 12561
rect -271 12527 -231 12561
rect -197 12527 -157 12561
rect -123 12527 -117 12561
rect -311 12489 -117 12527
rect -311 12455 -305 12489
rect -271 12455 -231 12489
rect -197 12455 -157 12489
rect -123 12455 -117 12489
rect -311 12417 -117 12455
rect 205 14462 743 14474
rect 205 14428 211 14462
rect 245 14428 293 14462
rect 327 14428 375 14462
rect 409 14428 457 14462
rect 491 14428 539 14462
rect 573 14428 621 14462
rect 655 14428 703 14462
rect 737 14428 743 14462
rect 205 14389 743 14428
rect 205 14355 211 14389
rect 245 14355 293 14389
rect 327 14355 375 14389
rect 409 14355 457 14389
rect 491 14355 539 14389
rect 573 14355 621 14389
rect 655 14355 703 14389
rect 737 14355 743 14389
rect 205 14316 743 14355
rect 205 14282 211 14316
rect 245 14282 293 14316
rect 327 14282 375 14316
rect 409 14282 457 14316
rect 491 14282 539 14316
rect 573 14282 621 14316
rect 655 14282 703 14316
rect 737 14282 743 14316
rect 205 14243 743 14282
rect 205 14209 211 14243
rect 245 14209 293 14243
rect 327 14209 375 14243
rect 409 14209 457 14243
rect 491 14209 539 14243
rect 573 14209 621 14243
rect 655 14209 703 14243
rect 737 14209 743 14243
rect 205 14170 743 14209
rect 205 14136 211 14170
rect 245 14136 293 14170
rect 327 14136 375 14170
rect 409 14136 457 14170
rect 491 14136 539 14170
rect 573 14136 621 14170
rect 655 14136 703 14170
rect 737 14136 743 14170
rect 205 14097 743 14136
rect 205 14063 211 14097
rect 245 14063 293 14097
rect 327 14063 375 14097
rect 409 14063 457 14097
rect 491 14063 539 14097
rect 573 14063 621 14097
rect 655 14063 703 14097
rect 737 14063 743 14097
rect 205 14029 743 14063
rect 205 14024 216 14029
rect 205 13990 211 14024
rect 205 13977 216 13990
rect 268 13977 281 14029
rect 333 13977 347 14029
rect 399 14024 413 14029
rect 465 14024 479 14029
rect 531 14024 545 14029
rect 409 13990 413 14024
rect 531 13990 539 14024
rect 399 13977 413 13990
rect 465 13977 479 13990
rect 531 13977 545 13990
rect 597 13977 611 14029
rect 663 13977 677 14029
rect 729 14024 743 14029
rect 737 13990 743 14024
rect 729 13977 743 13990
rect 205 13955 743 13977
rect 205 13951 216 13955
rect 205 13917 211 13951
rect 205 13903 216 13917
rect 268 13903 281 13955
rect 333 13903 347 13955
rect 399 13951 413 13955
rect 465 13951 479 13955
rect 531 13951 545 13955
rect 409 13917 413 13951
rect 531 13917 539 13951
rect 399 13903 413 13917
rect 465 13903 479 13917
rect 531 13903 545 13917
rect 597 13903 611 13955
rect 663 13903 677 13955
rect 729 13951 743 13955
rect 737 13917 743 13951
rect 729 13903 743 13917
rect 205 13881 743 13903
rect 205 13878 216 13881
rect 205 13844 211 13878
rect 205 13829 216 13844
rect 268 13829 281 13881
rect 333 13829 347 13881
rect 399 13878 413 13881
rect 465 13878 479 13881
rect 531 13878 545 13881
rect 409 13844 413 13878
rect 531 13844 539 13878
rect 399 13829 413 13844
rect 465 13829 479 13844
rect 531 13829 545 13844
rect 597 13829 611 13881
rect 663 13829 677 13881
rect 729 13878 743 13881
rect 737 13844 743 13878
rect 729 13829 743 13844
rect 205 13807 743 13829
rect 205 13805 216 13807
rect 205 13771 211 13805
rect 205 13755 216 13771
rect 268 13755 281 13807
rect 333 13755 347 13807
rect 399 13805 413 13807
rect 465 13805 479 13807
rect 531 13805 545 13807
rect 409 13771 413 13805
rect 531 13771 539 13805
rect 399 13755 413 13771
rect 465 13755 479 13771
rect 531 13755 545 13771
rect 597 13755 611 13807
rect 663 13755 677 13807
rect 729 13805 743 13807
rect 737 13771 743 13805
rect 729 13755 743 13771
rect 205 13733 743 13755
rect 205 13732 216 13733
rect 205 13698 211 13732
rect 205 13681 216 13698
rect 268 13681 281 13733
rect 333 13681 347 13733
rect 399 13732 413 13733
rect 465 13732 479 13733
rect 531 13732 545 13733
rect 409 13698 413 13732
rect 531 13698 539 13732
rect 399 13681 413 13698
rect 465 13681 479 13698
rect 531 13681 545 13698
rect 597 13681 611 13733
rect 663 13681 677 13733
rect 729 13732 743 13733
rect 737 13698 743 13732
rect 729 13681 743 13698
rect 205 13658 743 13681
rect 886 14029 1088 14035
rect 886 13977 887 14029
rect 939 13977 961 14029
rect 1013 13977 1035 14029
rect 1087 13977 1088 14029
rect 886 13955 1088 13977
rect 886 13903 887 13955
rect 939 13903 961 13955
rect 1013 13903 1035 13955
rect 1087 13903 1088 13955
rect 886 13881 1088 13903
rect 886 13829 887 13881
rect 939 13829 961 13881
rect 1013 13829 1035 13881
rect 1087 13829 1088 13881
rect 886 13807 1088 13829
rect 886 13755 887 13807
rect 939 13755 961 13807
rect 1013 13755 1035 13807
rect 1087 13755 1088 13807
rect 886 13733 1088 13755
rect 886 13681 887 13733
rect 939 13681 961 13733
rect 1013 13681 1035 13733
rect 1087 13681 1088 13733
rect 886 13675 1088 13681
rect 205 13624 211 13658
rect 245 13624 293 13658
rect 327 13624 375 13658
rect 409 13624 457 13658
rect 491 13624 539 13658
rect 573 13624 621 13658
rect 655 13624 703 13658
rect 737 13624 743 13658
rect 205 13584 743 13624
rect 205 13550 211 13584
rect 245 13550 293 13584
rect 327 13550 375 13584
rect 409 13550 457 13584
rect 491 13550 539 13584
rect 573 13550 621 13584
rect 655 13550 703 13584
rect 737 13550 743 13584
rect 205 13510 743 13550
rect 205 13476 211 13510
rect 245 13476 293 13510
rect 327 13476 375 13510
rect 409 13476 457 13510
rect 491 13476 539 13510
rect 573 13476 621 13510
rect 655 13476 703 13510
rect 737 13476 743 13510
rect 205 13436 743 13476
rect 205 13402 211 13436
rect 245 13402 293 13436
rect 327 13402 375 13436
rect 409 13402 457 13436
rect 491 13402 539 13436
rect 573 13402 621 13436
rect 655 13402 703 13436
rect 737 13402 743 13436
rect 205 13362 743 13402
rect 205 13328 211 13362
rect 245 13328 293 13362
rect 327 13328 375 13362
rect 409 13328 457 13362
rect 491 13328 539 13362
rect 573 13328 621 13362
rect 655 13328 703 13362
rect 737 13328 743 13362
rect 205 13288 743 13328
rect 205 13254 211 13288
rect 245 13254 293 13288
rect 327 13254 375 13288
rect 409 13254 457 13288
rect 491 13254 539 13288
rect 573 13254 621 13288
rect 655 13254 703 13288
rect 737 13254 743 13288
rect 205 13214 743 13254
rect 205 13180 211 13214
rect 245 13180 293 13214
rect 327 13180 375 13214
rect 409 13180 457 13214
rect 491 13180 539 13214
rect 573 13180 621 13214
rect 655 13180 703 13214
rect 737 13180 743 13214
rect 205 13140 743 13180
rect 205 13106 211 13140
rect 245 13106 293 13140
rect 327 13106 375 13140
rect 409 13106 457 13140
rect 491 13106 539 13140
rect 573 13106 621 13140
rect 655 13106 703 13140
rect 737 13106 743 13140
rect 205 13066 743 13106
rect 205 13032 211 13066
rect 245 13032 293 13066
rect 327 13032 375 13066
rect 409 13032 457 13066
rect 491 13032 539 13066
rect 573 13032 621 13066
rect 655 13032 703 13066
rect 737 13032 743 13066
rect 205 12992 743 13032
rect 205 12958 211 12992
rect 245 12958 293 12992
rect 327 12958 375 12992
rect 409 12958 457 12992
rect 491 12958 539 12992
rect 573 12958 621 12992
rect 655 12958 703 12992
rect 737 12958 743 12992
rect 205 12918 743 12958
rect 205 12884 211 12918
rect 245 12884 293 12918
rect 327 12884 375 12918
rect 409 12884 457 12918
rect 491 12884 539 12918
rect 573 12884 621 12918
rect 655 12884 703 12918
rect 737 12884 743 12918
rect 205 12844 743 12884
rect 205 12810 211 12844
rect 245 12810 293 12844
rect 327 12810 375 12844
rect 409 12810 457 12844
rect 491 12810 539 12844
rect 573 12810 621 12844
rect 655 12810 703 12844
rect 737 12810 743 12844
rect 205 12770 743 12810
rect 205 12736 211 12770
rect 245 12736 293 12770
rect 327 12736 375 12770
rect 409 12736 457 12770
rect 491 12736 539 12770
rect 573 12736 621 12770
rect 655 12736 703 12770
rect 737 12736 743 12770
rect 205 12696 743 12736
rect 205 12662 211 12696
rect 245 12662 293 12696
rect 327 12662 375 12696
rect 409 12662 457 12696
rect 491 12662 539 12696
rect 573 12662 621 12696
rect 655 12662 703 12696
rect 737 12662 743 12696
rect 205 12622 743 12662
rect 205 12588 211 12622
rect 245 12588 293 12622
rect 327 12588 375 12622
rect 409 12588 457 12622
rect 491 12588 539 12622
rect 573 12588 621 12622
rect 655 12588 703 12622
rect 737 12588 743 12622
rect 205 12548 743 12588
rect 205 12514 211 12548
rect 245 12514 293 12548
rect 327 12514 375 12548
rect 409 12514 457 12548
rect 491 12514 539 12548
rect 573 12514 621 12548
rect 655 12514 703 12548
rect 737 12514 743 12548
rect 205 12474 743 12514
rect 205 12440 211 12474
rect 245 12440 293 12474
rect 327 12440 375 12474
rect 409 12440 457 12474
rect 491 12440 539 12474
rect 573 12440 621 12474
rect 655 12440 703 12474
rect 737 12440 743 12474
rect 205 12428 743 12440
rect -311 12383 -305 12417
rect -271 12383 -231 12417
rect -197 12383 -157 12417
rect -123 12383 -117 12417
rect -311 12345 -117 12383
rect -311 12311 -305 12345
rect -271 12311 -231 12345
rect -197 12311 -157 12345
rect -123 12311 -117 12345
rect -311 12273 -117 12311
rect -311 12239 -305 12273
rect -271 12239 -231 12273
rect -197 12239 -157 12273
rect -123 12239 -117 12273
rect -311 12201 -117 12239
rect -311 12167 -305 12201
rect -271 12167 -231 12201
rect -197 12167 -157 12201
rect -123 12167 -117 12201
rect -311 12166 -117 12167
rect -311 12095 -305 12166
rect -253 12114 -240 12166
rect -188 12114 -175 12166
rect -271 12095 -231 12114
rect -197 12095 -157 12114
rect -123 12095 -117 12166
rect -68 12114 -62 12166
rect -10 12114 8 12166
rect 60 12114 78 12166
rect 130 12114 148 12166
rect 200 12114 218 12166
rect 270 12114 289 12166
rect 341 12114 347 12166
tri 347 12114 353 12120 nw
rect -311 12057 -117 12095
rect -311 12023 -305 12057
rect -271 12023 -231 12057
rect -197 12023 -157 12057
rect -123 12023 -117 12057
rect -311 11985 -117 12023
rect -311 11951 -305 11985
rect -271 11951 -231 11985
rect -197 11951 -157 11985
rect -123 11951 -117 11985
rect -311 11913 -117 11951
rect -311 11879 -305 11913
rect -271 11879 -231 11913
rect -197 11879 -157 11913
rect -123 11879 -117 11913
rect -311 11841 -117 11879
rect -311 11807 -305 11841
rect -271 11807 -231 11841
rect -197 11807 -157 11841
rect -123 11807 -117 11841
rect -311 11769 -117 11807
rect -311 11735 -305 11769
rect -271 11735 -231 11769
rect -197 11735 -157 11769
rect -123 11735 -117 11769
rect -311 11697 -117 11735
rect -311 11663 -305 11697
rect -271 11663 -231 11697
rect -197 11663 -157 11697
rect -123 11663 -117 11697
rect -311 11625 -117 11663
rect -311 11591 -305 11625
rect -271 11591 -231 11625
rect -197 11591 -157 11625
rect -123 11591 -117 11625
rect -311 11553 -117 11591
rect -311 11519 -305 11553
rect -271 11519 -231 11553
rect -197 11519 -157 11553
rect -123 11519 -117 11553
rect -311 11481 -117 11519
rect -311 11447 -305 11481
rect -271 11447 -231 11481
rect -197 11447 -157 11481
rect -123 11447 -117 11481
rect -311 11409 -117 11447
rect -311 11375 -305 11409
rect -271 11375 -231 11409
rect -197 11375 -157 11409
rect -123 11375 -117 11409
rect -311 11337 -117 11375
rect -311 11303 -305 11337
rect -271 11303 -231 11337
rect -197 11303 -157 11337
rect -123 11303 -117 11337
rect -311 11265 -117 11303
rect -311 11231 -305 11265
rect -271 11231 -231 11265
rect -197 11231 -157 11265
rect -123 11231 -117 11265
rect -311 11193 -117 11231
rect -311 11159 -305 11193
rect -271 11159 -231 11193
rect -197 11159 -157 11193
rect -123 11159 -117 11193
rect -311 11121 -117 11159
rect -311 11087 -305 11121
rect -271 11087 -231 11121
rect -197 11087 -157 11121
rect -123 11087 -117 11121
rect -311 11049 -117 11087
rect -311 11015 -305 11049
rect -271 11015 -231 11049
rect -197 11015 -157 11049
rect -123 11015 -117 11049
rect -311 10977 -117 11015
rect -311 10943 -305 10977
rect -271 10943 -231 10977
rect -197 10943 -157 10977
rect -123 10943 -117 10977
rect -311 10905 -117 10943
rect -311 10871 -305 10905
rect -271 10871 -231 10905
rect -197 10871 -157 10905
rect -123 10871 -117 10905
rect -311 10833 -117 10871
rect -311 10799 -305 10833
rect -271 10799 -231 10833
rect -197 10799 -157 10833
rect -123 10799 -117 10833
rect -311 10761 -117 10799
rect -311 10727 -305 10761
rect -271 10727 -231 10761
rect -197 10727 -157 10761
rect -123 10727 -117 10761
rect -311 10689 -117 10727
rect -311 10655 -305 10689
rect -271 10655 -231 10689
rect -197 10655 -157 10689
rect -123 10655 -117 10689
rect -311 10617 -117 10655
rect -311 10583 -305 10617
rect -271 10583 -231 10617
rect -197 10583 -157 10617
rect -123 10583 -117 10617
rect -311 10545 -117 10583
rect -311 10511 -305 10545
rect -271 10511 -231 10545
rect -197 10511 -157 10545
rect -123 10511 -117 10545
rect -311 10473 -117 10511
rect -311 10439 -305 10473
rect -271 10439 -231 10473
rect -197 10439 -157 10473
rect -123 10439 -117 10473
rect -311 10401 -117 10439
rect -311 10367 -305 10401
rect -271 10367 -231 10401
rect -197 10367 -157 10401
rect -123 10367 -117 10401
rect -311 10329 -117 10367
rect -311 10295 -305 10329
rect -271 10295 -231 10329
rect -197 10295 -157 10329
rect -123 10295 -117 10329
rect -311 10257 -117 10295
rect -311 10223 -305 10257
rect -271 10223 -231 10257
rect -197 10223 -157 10257
rect -123 10223 -117 10257
rect -311 10185 -117 10223
rect -311 10151 -305 10185
rect -271 10151 -231 10185
rect -197 10151 -157 10185
rect -123 10151 -117 10185
rect -311 10113 -117 10151
rect -311 10079 -305 10113
rect -271 10079 -231 10113
rect -197 10079 -157 10113
rect -123 10079 -117 10113
rect -311 10041 -117 10079
rect -311 10007 -305 10041
rect -271 10007 -231 10041
rect -197 10007 -157 10041
rect -123 10007 -117 10041
rect -311 9969 -117 10007
rect -311 9935 -305 9969
rect -271 9935 -231 9969
rect -197 9935 -157 9969
rect -123 9935 -117 9969
rect -311 9897 -117 9935
rect -311 9863 -305 9897
rect -271 9863 -231 9897
rect -197 9863 -157 9897
rect -123 9863 -117 9897
rect -311 9825 -117 9863
rect -311 9791 -305 9825
rect -271 9791 -231 9825
rect -197 9791 -157 9825
rect -123 9791 -117 9825
rect -311 9753 -117 9791
rect -311 9719 -305 9753
rect -271 9719 -231 9753
rect -197 9719 -157 9753
rect -123 9719 -117 9753
rect -311 9681 -117 9719
rect -311 9647 -305 9681
rect -271 9647 -231 9681
rect -197 9647 -157 9681
rect -123 9647 -117 9681
rect -311 9609 -117 9647
rect -311 9575 -305 9609
rect -271 9575 -231 9609
rect -197 9575 -157 9609
rect -123 9575 -117 9609
rect -311 9537 -117 9575
rect -311 9503 -305 9537
rect -271 9503 -231 9537
rect -197 9503 -157 9537
rect -123 9503 -117 9537
rect -311 9465 -117 9503
rect -311 9431 -305 9465
rect -271 9431 -231 9465
rect -197 9431 -157 9465
rect -123 9431 -117 9465
rect -311 9393 -117 9431
rect -311 9359 -305 9393
rect -271 9359 -231 9393
rect -197 9359 -157 9393
rect -123 9359 -117 9393
rect -311 9321 -117 9359
rect -311 9287 -305 9321
rect -271 9287 -231 9321
rect -197 9287 -157 9321
rect -123 9287 -117 9321
rect -311 9249 -117 9287
rect -311 9215 -305 9249
rect -271 9215 -231 9249
rect -197 9215 -157 9249
rect -123 9215 -117 9249
rect -311 9177 -117 9215
rect -311 9143 -305 9177
rect -271 9143 -231 9177
rect -197 9143 -157 9177
rect -123 9143 -117 9177
rect -311 9105 -117 9143
rect -311 9071 -305 9105
rect -271 9071 -231 9105
rect -197 9071 -157 9105
rect -123 9071 -117 9105
rect -311 9033 -117 9071
rect -311 8999 -305 9033
rect -271 8999 -231 9033
rect -197 8999 -157 9033
rect -123 8999 -117 9033
rect -311 8961 -117 8999
rect -311 8927 -305 8961
rect -271 8927 -231 8961
rect -197 8927 -157 8961
rect -123 8927 -117 8961
rect -311 8889 -117 8927
rect -311 8855 -305 8889
rect -271 8855 -231 8889
rect -197 8855 -157 8889
rect -123 8855 -117 8889
rect -311 8817 -117 8855
rect -311 8783 -305 8817
rect -271 8783 -231 8817
rect -197 8783 -157 8817
rect -123 8783 -117 8817
rect -311 8745 -117 8783
rect -311 8711 -305 8745
rect -271 8711 -231 8745
rect -197 8711 -157 8745
rect -123 8711 -117 8745
rect -311 8673 -117 8711
rect -311 8639 -305 8673
rect -271 8639 -231 8673
rect -197 8639 -157 8673
rect -123 8639 -117 8673
rect -311 8601 -117 8639
rect -311 8567 -305 8601
rect -271 8567 -231 8601
rect -197 8567 -157 8601
rect -123 8567 -117 8601
rect -311 8529 -117 8567
rect -311 8495 -305 8529
rect -271 8495 -231 8529
rect -197 8495 -157 8529
rect -123 8495 -117 8529
rect -311 8457 -117 8495
rect -311 8423 -305 8457
rect -271 8423 -231 8457
rect -197 8423 -157 8457
rect -123 8423 -117 8457
rect -311 8385 -117 8423
rect -311 8351 -305 8385
rect -271 8351 -231 8385
rect -197 8351 -157 8385
rect -123 8351 -117 8385
rect -311 8313 -117 8351
rect -311 8279 -305 8313
rect -271 8279 -231 8313
rect -197 8279 -157 8313
rect -123 8279 -117 8313
rect -311 8241 -117 8279
rect -311 8207 -305 8241
rect -271 8207 -231 8241
rect -197 8207 -157 8241
rect -123 8207 -117 8241
rect -311 8168 -117 8207
rect -311 8134 -305 8168
rect -271 8134 -231 8168
rect -197 8134 -157 8168
rect -123 8134 -117 8168
rect -311 8095 -117 8134
rect -311 8061 -305 8095
rect -271 8061 -231 8095
rect -197 8061 -157 8095
rect -123 8061 -117 8095
rect -311 8022 -117 8061
rect -311 7988 -305 8022
rect -271 7988 -231 8022
rect -197 7988 -157 8022
rect -123 7988 -117 8022
rect -311 7949 -117 7988
rect -311 7915 -305 7949
rect -271 7915 -231 7949
rect -197 7915 -157 7949
rect -123 7915 -117 7949
rect -311 7876 -117 7915
rect -311 7842 -305 7876
rect -271 7842 -231 7876
rect -197 7842 -157 7876
rect -123 7842 -117 7876
rect -311 7803 -117 7842
rect -311 7769 -305 7803
rect -271 7769 -231 7803
rect -197 7769 -157 7803
rect -123 7769 -117 7803
rect -311 7730 -117 7769
rect -311 7696 -305 7730
rect -271 7696 -231 7730
rect -197 7696 -157 7730
rect -123 7696 -117 7730
rect -311 7657 -117 7696
rect -311 7623 -305 7657
rect -271 7623 -231 7657
rect -197 7623 -157 7657
rect -123 7623 -117 7657
rect -311 7584 -117 7623
rect -311 7550 -305 7584
rect -271 7550 -231 7584
rect -197 7550 -157 7584
rect -123 7550 -117 7584
rect -311 7511 -117 7550
rect -311 7477 -305 7511
rect -271 7477 -231 7511
rect -197 7477 -157 7511
rect -123 7477 -117 7511
rect -311 7438 -117 7477
rect -311 7404 -305 7438
rect -271 7404 -231 7438
rect -197 7404 -157 7438
rect -123 7404 -117 7438
rect -311 7365 -117 7404
rect -311 7331 -305 7365
rect -271 7331 -231 7365
rect -197 7331 -157 7365
rect -123 7331 -117 7365
rect -311 7292 -117 7331
rect -311 7258 -305 7292
rect -271 7258 -231 7292
rect -197 7258 -157 7292
rect -123 7258 -117 7292
rect -311 7219 -117 7258
rect -311 7185 -305 7219
rect -271 7185 -231 7219
rect -197 7185 -157 7219
rect -123 7185 -117 7219
rect -311 7146 -117 7185
rect -311 7112 -305 7146
rect -271 7112 -231 7146
rect -197 7112 -157 7146
rect -123 7112 -117 7146
rect -311 7073 -117 7112
rect -311 7039 -305 7073
rect -271 7039 -231 7073
rect -197 7039 -157 7073
rect -123 7039 -117 7073
rect -311 7000 -117 7039
rect -311 6966 -305 7000
rect -271 6966 -231 7000
rect -197 6966 -157 7000
rect -123 6966 -117 7000
rect -311 6927 -117 6966
rect -311 6893 -305 6927
rect -271 6893 -231 6927
rect -197 6893 -157 6927
rect -123 6893 -117 6927
rect -311 6854 -117 6893
rect -311 6820 -305 6854
rect -271 6820 -231 6854
rect -197 6820 -157 6854
rect -123 6820 -117 6854
rect -311 6781 -117 6820
rect -311 6747 -305 6781
rect -271 6747 -231 6781
rect -197 6747 -157 6781
rect -123 6747 -117 6781
rect -311 6708 -117 6747
rect -311 6674 -305 6708
rect -271 6674 -231 6708
rect -197 6674 -157 6708
rect -123 6674 -117 6708
rect -311 6635 -117 6674
rect -311 6601 -305 6635
rect -271 6601 -231 6635
rect -197 6601 -157 6635
rect -123 6601 -117 6635
rect -311 6562 -117 6601
rect -311 6528 -305 6562
rect -271 6528 -231 6562
rect -197 6528 -157 6562
rect -123 6528 -117 6562
rect -311 6489 -117 6528
rect -311 6455 -305 6489
rect -271 6455 -231 6489
rect -197 6455 -157 6489
rect -123 6455 -117 6489
rect -311 6416 -117 6455
rect -311 6391 -305 6416
rect -271 6391 -231 6416
rect -197 6391 -157 6416
rect -123 6391 -117 6416
tri -22 6397 -16 6403 sw
rect -311 6339 -310 6391
rect -258 6339 -240 6391
rect -188 6339 -170 6391
rect -118 6339 -117 6391
rect -311 6321 -305 6339
rect -271 6321 -231 6339
rect -197 6321 -157 6339
rect -123 6321 -117 6339
rect -311 6269 -310 6321
rect -258 6269 -240 6321
rect -188 6269 -170 6321
rect -118 6269 -117 6321
rect -311 6251 -305 6269
rect -271 6251 -231 6269
rect -197 6251 -157 6269
rect -123 6251 -117 6269
rect -311 6199 -310 6251
rect -258 6199 -240 6251
rect -188 6199 -170 6251
rect -118 6199 -117 6251
rect -311 6197 -117 6199
rect -311 6181 -305 6197
rect -271 6181 -231 6197
rect -197 6181 -157 6197
rect -123 6181 -117 6197
rect -311 6129 -310 6181
rect -258 6129 -240 6181
rect -188 6129 -170 6181
rect -118 6129 -117 6181
rect -311 6124 -117 6129
rect -311 6111 -305 6124
rect -271 6111 -231 6124
rect -197 6111 -157 6124
rect -123 6111 -117 6124
rect -311 6059 -310 6111
rect -258 6059 -240 6111
rect -188 6059 -170 6111
rect -118 6059 -117 6111
rect -311 6051 -117 6059
rect -311 6041 -305 6051
rect -271 6041 -231 6051
rect -197 6041 -157 6051
rect -123 6041 -117 6051
rect -311 5989 -310 6041
rect -258 5989 -240 6041
rect -188 5989 -170 6041
rect -118 5989 -117 6041
rect -311 5978 -117 5989
rect -311 5971 -305 5978
rect -271 5971 -231 5978
rect -197 5971 -157 5978
rect -123 5971 -117 5978
rect -311 5919 -310 5971
rect -258 5919 -240 5971
rect -188 5919 -170 5971
rect -118 5919 -117 5971
rect -311 5905 -117 5919
rect -311 5901 -305 5905
rect -271 5901 -231 5905
rect -197 5901 -157 5905
rect -123 5901 -117 5905
rect -311 5849 -310 5901
rect -258 5849 -240 5901
rect -188 5849 -170 5901
rect -118 5849 -117 5901
rect -311 5832 -117 5849
rect -311 5830 -305 5832
rect -271 5830 -231 5832
rect -197 5830 -157 5832
rect -123 5830 -117 5832
rect -311 5778 -310 5830
rect -258 5778 -240 5830
rect -188 5778 -170 5830
rect -118 5778 -117 5830
rect -311 5759 -117 5778
rect -68 6391 -16 6397
rect -68 6321 -16 6339
rect -68 6251 -16 6269
rect -68 6181 -16 6199
rect -68 6111 -16 6129
rect -68 6041 -16 6059
rect -68 5971 -16 5989
rect -68 5901 -16 5919
rect -68 5830 -16 5849
rect -68 5772 -16 5778
tri -22 5766 -16 5772 nw
rect -311 5725 -305 5759
rect -271 5725 -231 5759
rect -197 5725 -157 5759
rect -123 5725 -117 5759
rect -311 5686 -117 5725
rect -311 5652 -305 5686
rect -271 5652 -231 5686
rect -197 5652 -157 5686
rect -123 5652 -117 5686
rect -311 5613 -117 5652
rect -311 5579 -305 5613
rect -271 5579 -231 5613
rect -197 5579 -157 5613
rect -123 5579 -117 5613
rect -311 5540 -117 5579
rect -311 5506 -305 5540
rect -271 5506 -231 5540
rect -197 5506 -157 5540
rect -123 5506 -117 5540
rect -311 5467 -117 5506
rect -311 5433 -305 5467
rect -271 5433 -231 5467
rect -197 5433 -157 5467
rect -123 5433 -117 5467
rect -311 5394 -117 5433
rect -311 5360 -305 5394
rect -271 5360 -231 5394
rect -197 5360 -157 5394
rect -123 5360 -117 5394
rect -311 5321 -117 5360
rect -311 5287 -305 5321
rect -271 5287 -231 5321
rect -197 5287 -157 5321
rect -123 5287 -117 5321
rect -311 5248 -117 5287
rect -311 5214 -305 5248
rect -271 5214 -231 5248
rect -197 5214 -157 5248
rect -123 5214 -117 5248
rect -311 5175 -117 5214
rect -311 5141 -305 5175
rect -271 5141 -231 5175
rect -197 5141 -157 5175
rect -123 5141 -117 5175
rect -311 5102 -117 5141
rect -311 5070 -305 5102
rect -271 5070 -231 5102
rect -197 5070 -157 5102
rect -123 5070 -117 5102
tri -22 5076 -16 5082 sw
rect -311 5018 -310 5070
rect -258 5018 -240 5070
rect -188 5018 -170 5070
rect -118 5018 -117 5070
rect -311 5004 -305 5018
rect -271 5004 -231 5018
rect -197 5004 -157 5018
rect -123 5004 -117 5018
rect -311 4952 -310 5004
rect -258 4952 -240 5004
rect -188 4952 -170 5004
rect -118 4952 -117 5004
rect -311 4938 -305 4952
rect -271 4938 -231 4952
rect -197 4938 -157 4952
rect -123 4938 -117 4952
rect -311 4886 -310 4938
rect -258 4886 -240 4938
rect -188 4886 -170 4938
rect -118 4886 -117 4938
rect -311 4883 -117 4886
rect -311 4872 -305 4883
rect -271 4872 -231 4883
rect -197 4872 -157 4883
rect -123 4872 -117 4883
rect -311 4820 -310 4872
rect -258 4820 -240 4872
rect -188 4820 -170 4872
rect -118 4820 -117 4872
rect -311 4810 -117 4820
rect -311 4806 -305 4810
rect -271 4806 -231 4810
rect -197 4806 -157 4810
rect -123 4806 -117 4810
rect -311 4754 -310 4806
rect -258 4754 -240 4806
rect -188 4754 -170 4806
rect -118 4754 -117 4806
rect -311 4740 -117 4754
rect -311 4688 -310 4740
rect -258 4688 -240 4740
rect -188 4688 -170 4740
rect -118 4688 -117 4740
rect -311 4674 -117 4688
rect -311 4622 -310 4674
rect -258 4622 -240 4674
rect -188 4622 -170 4674
rect -118 4622 -117 4674
rect -311 4607 -117 4622
rect -311 4555 -310 4607
rect -258 4555 -240 4607
rect -188 4555 -170 4607
rect -118 4555 -117 4607
rect -311 4540 -117 4555
rect -311 4488 -310 4540
rect -258 4488 -240 4540
rect -188 4488 -170 4540
rect -118 4488 -117 4540
rect -311 4484 -305 4488
rect -271 4484 -231 4488
rect -197 4484 -157 4488
rect -123 4484 -117 4488
rect -311 4473 -117 4484
rect -311 4421 -310 4473
rect -258 4421 -240 4473
rect -188 4421 -170 4473
rect -118 4421 -117 4473
rect -311 4411 -305 4421
rect -271 4411 -231 4421
rect -197 4411 -157 4421
rect -123 4411 -117 4421
rect -311 4406 -117 4411
rect -311 4354 -310 4406
rect -258 4354 -240 4406
rect -188 4354 -170 4406
rect -118 4354 -117 4406
rect -311 4339 -305 4354
rect -271 4339 -231 4354
rect -197 4339 -157 4354
rect -123 4339 -117 4354
rect -311 4287 -310 4339
rect -258 4287 -240 4339
rect -188 4287 -170 4339
rect -118 4287 -117 4339
rect -311 4272 -305 4287
rect -271 4272 -231 4287
rect -197 4272 -157 4287
rect -123 4272 -117 4287
rect -311 4220 -310 4272
rect -258 4220 -240 4272
rect -188 4220 -170 4272
rect -118 4220 -117 4272
rect -311 4205 -305 4220
rect -271 4205 -231 4220
rect -197 4205 -157 4220
rect -123 4205 -117 4220
rect -311 4153 -310 4205
rect -258 4153 -240 4205
rect -188 4153 -170 4205
rect -118 4153 -117 4205
rect -311 4138 -305 4153
rect -271 4138 -231 4153
rect -197 4138 -157 4153
rect -123 4138 -117 4153
rect -311 4086 -310 4138
rect -258 4086 -240 4138
rect -188 4086 -170 4138
rect -118 4086 -117 4138
rect -311 4080 -117 4086
rect -311 4071 -305 4080
rect -271 4071 -231 4080
rect -197 4071 -157 4080
rect -123 4071 -117 4080
rect -311 4019 -310 4071
rect -258 4019 -240 4071
rect -188 4019 -170 4071
rect -118 4019 -117 4071
rect -311 4007 -117 4019
rect -311 3973 -305 4007
rect -271 3973 -231 4007
rect -197 3973 -157 4007
rect -123 3973 -117 4007
rect -311 3934 -117 3973
rect -311 3900 -305 3934
rect -271 3900 -231 3934
rect -197 3900 -157 3934
rect -123 3900 -117 3934
rect -311 3861 -117 3900
rect -311 3827 -305 3861
rect -271 3827 -231 3861
rect -197 3827 -157 3861
rect -123 3827 -117 3861
rect -311 3788 -117 3827
rect -311 3754 -305 3788
rect -271 3754 -231 3788
rect -197 3754 -157 3788
rect -123 3754 -117 3788
rect -311 3715 -117 3754
rect -311 3681 -305 3715
rect -271 3681 -231 3715
rect -197 3681 -157 3715
rect -123 3681 -117 3715
rect -311 3642 -117 3681
rect -311 3608 -305 3642
rect -271 3608 -231 3642
rect -197 3608 -157 3642
rect -123 3608 -117 3642
rect -311 3569 -117 3608
rect -311 3535 -305 3569
rect -271 3535 -231 3569
rect -197 3535 -157 3569
rect -123 3535 -117 3569
rect -311 3496 -117 3535
rect -311 3462 -305 3496
rect -271 3462 -231 3496
rect -197 3462 -157 3496
rect -123 3462 -117 3496
rect -311 3450 -117 3462
rect -68 5070 -16 5076
rect -68 5016 -16 5018
rect -68 5010 936 5016
rect -68 5004 28 5010
rect -16 4976 28 5004
rect 62 4976 106 5010
rect 140 4976 184 5010
rect 218 4976 262 5010
rect 296 4976 340 5010
rect 374 4976 418 5010
rect 452 4976 496 5010
rect 530 4976 574 5010
rect 608 4976 652 5010
rect 686 4976 730 5010
rect 764 4976 808 5010
rect 842 4976 936 5010
rect -16 4970 936 4976
rect -68 4940 -62 4952
rect -28 4940 -16 4952
rect -68 4938 -16 4940
tri -16 4939 15 4970 nw
tri 808 4939 839 4970 ne
rect 839 4939 936 4970
tri 839 4933 845 4939 ne
rect 845 4933 936 4939
rect -68 4872 -62 4886
rect -28 4872 -16 4886
tri 845 4870 908 4933 ne
rect 908 4870 936 4933
rect -68 4806 -62 4820
rect -28 4806 -16 4820
rect -68 4740 -62 4754
rect -28 4740 -16 4754
rect -68 4682 -16 4688
rect -68 4674 -62 4682
rect -28 4674 -16 4682
rect -68 4609 -16 4622
rect -68 4607 -62 4609
rect -28 4607 -16 4609
rect -68 4540 -16 4555
rect -68 4473 -16 4488
rect -68 4406 -16 4421
rect -68 4339 -16 4354
rect -68 4283 -62 4287
rect -28 4283 -16 4287
rect -68 4272 -16 4283
rect -68 4210 -62 4220
rect -28 4210 -16 4220
rect -68 4205 -16 4210
rect -68 4138 -62 4153
rect -28 4138 -16 4153
rect -68 4071 -62 4086
rect -28 4071 -16 4086
rect -68 3992 -62 4019
rect -28 4013 -16 4019
rect -28 3992 -22 4013
tri -22 4007 -16 4013 nw
rect 153 4842 703 4860
rect 153 4808 231 4842
rect 265 4808 303 4842
rect 337 4808 375 4842
rect 409 4808 447 4842
rect 481 4808 519 4842
rect 553 4808 703 4842
rect 153 4790 703 4808
rect 153 4782 249 4790
tri 249 4782 257 4790 nw
tri 599 4782 607 4790 ne
rect 607 4782 703 4790
rect 153 4778 223 4782
rect 153 4744 171 4778
rect 205 4744 223 4778
tri 223 4756 249 4782 nw
tri 607 4756 633 4782 ne
rect 153 4702 223 4744
rect 153 4691 171 4702
rect 205 4691 223 4702
rect 153 4639 162 4691
rect 214 4639 223 4691
rect 633 4748 651 4782
rect 685 4748 703 4782
rect 633 4708 703 4748
rect 633 4674 651 4708
rect 685 4674 703 4708
rect 153 4626 223 4639
rect 153 4625 171 4626
rect 205 4625 223 4626
rect 153 4573 162 4625
rect 214 4573 223 4625
rect 153 4558 223 4573
rect 153 4506 162 4558
rect 214 4506 223 4558
rect 153 4491 223 4506
rect 153 4439 162 4491
rect 214 4439 223 4491
rect 153 4424 223 4439
rect 153 4372 162 4424
rect 214 4372 223 4424
rect 153 4364 171 4372
rect 205 4364 223 4372
rect 153 4357 223 4364
rect 153 4305 162 4357
rect 214 4305 223 4357
rect 153 4290 171 4305
rect 205 4290 223 4305
rect 153 4238 162 4290
rect 214 4238 223 4290
rect 153 4223 171 4238
rect 205 4223 223 4238
rect 153 4171 162 4223
rect 214 4171 223 4223
rect 153 4170 223 4171
rect 153 4136 171 4170
rect 205 4136 223 4170
rect 153 4093 223 4136
rect 153 4059 171 4093
rect 205 4059 223 4093
rect 153 4016 223 4059
rect -68 3954 -22 3992
rect -68 3920 -62 3954
rect -28 3920 -22 3954
rect -68 3882 -22 3920
rect -68 3848 -62 3882
rect -28 3848 -22 3882
rect -68 3810 -22 3848
rect -68 3776 -62 3810
rect -28 3776 -22 3810
rect -68 3738 -22 3776
rect -68 3704 -62 3738
rect -28 3704 -22 3738
rect -68 3666 -22 3704
rect -68 3632 -62 3666
rect -28 3632 -22 3666
rect -68 3594 -22 3632
rect -68 3560 -62 3594
rect -28 3560 -22 3594
rect 153 3982 171 4016
rect 205 3982 223 4016
rect 153 3939 223 3982
rect 153 3905 171 3939
rect 205 3905 223 3939
rect 153 3862 223 3905
rect 153 3828 171 3862
rect 205 3828 223 3862
rect 153 3785 223 3828
rect 153 3751 171 3785
rect 205 3751 223 3785
rect 278 4658 579 4670
rect 278 4624 284 4658
rect 318 4624 539 4658
rect 573 4624 579 4658
rect 278 4583 579 4624
rect 278 4549 284 4583
rect 318 4549 539 4583
rect 573 4549 579 4583
rect 278 4508 579 4549
rect 278 4474 284 4508
rect 318 4474 539 4508
rect 573 4474 579 4508
rect 278 4433 579 4474
rect 278 4399 284 4433
rect 318 4399 539 4433
rect 573 4399 579 4433
rect 278 4357 579 4399
rect 278 4323 284 4357
rect 318 4323 539 4357
rect 573 4323 579 4357
rect 278 4281 579 4323
rect 278 4247 284 4281
rect 318 4247 539 4281
rect 573 4247 579 4281
rect 278 4205 579 4247
rect 278 4171 284 4205
rect 318 4171 539 4205
rect 573 4171 579 4205
rect 278 4129 579 4171
rect 278 4095 284 4129
rect 318 4095 539 4129
rect 573 4095 579 4129
rect 278 4053 579 4095
rect 278 4019 284 4053
rect 318 4019 539 4053
rect 573 4019 579 4053
rect 278 3977 579 4019
rect 278 3943 284 3977
rect 318 3943 539 3977
rect 573 3943 579 3977
rect 278 3901 579 3943
rect 278 3867 284 3901
rect 318 3867 539 3901
rect 573 3867 579 3901
rect 278 3825 579 3867
rect 278 3791 284 3825
rect 318 3791 539 3825
rect 573 3791 579 3825
rect 278 3779 579 3791
rect 633 4634 703 4674
rect 633 4600 651 4634
rect 685 4600 703 4634
rect 633 4561 703 4600
rect 633 4527 651 4561
rect 685 4527 703 4561
rect 633 4488 703 4527
rect 633 4454 651 4488
rect 685 4454 703 4488
rect 633 4415 703 4454
rect 633 4381 651 4415
rect 685 4381 703 4415
rect 633 4342 703 4381
rect 633 4308 651 4342
rect 685 4308 703 4342
rect 633 4269 703 4308
rect 633 4235 651 4269
rect 685 4235 703 4269
rect 633 4196 703 4235
rect 633 4162 651 4196
rect 685 4162 703 4196
rect 633 4123 703 4162
rect 633 4089 651 4123
rect 685 4089 703 4123
rect 633 4050 703 4089
rect 633 4016 651 4050
rect 685 4016 703 4050
rect 633 3977 703 4016
rect 633 3943 651 3977
rect 685 3943 703 3977
rect 633 3904 703 3943
rect 633 3870 651 3904
rect 685 3870 703 3904
rect 633 3831 703 3870
rect 633 3797 651 3831
rect 685 3797 703 3831
rect 153 3708 223 3751
rect 153 3674 171 3708
rect 205 3674 223 3708
rect 633 3758 703 3797
rect 633 3724 651 3758
rect 685 3724 703 3758
rect 153 3631 223 3674
rect 364 3694 410 3706
rect 364 3660 370 3694
rect 404 3660 410 3694
rect 633 3685 703 3724
rect 153 3597 171 3631
rect 205 3625 223 3631
tri 223 3625 231 3633 sw
rect 205 3621 231 3625
tri 231 3621 235 3625 sw
rect 364 3621 410 3660
rect 205 3597 235 3621
rect 153 3587 235 3597
tri 235 3587 269 3621 sw
rect 364 3587 370 3621
rect 404 3587 410 3621
rect 153 3586 269 3587
tri 269 3586 270 3587 sw
rect 153 3585 270 3586
tri 270 3585 271 3586 sw
rect 153 3563 271 3585
tri 271 3563 293 3585 sw
tri 153 3561 155 3563 ne
rect 155 3561 293 3563
tri 293 3561 295 3563 sw
rect -68 3522 -22 3560
tri 155 3555 161 3561 ne
rect -68 3488 -62 3522
rect -28 3488 -22 3522
rect -68 3450 -22 3488
rect -824 3395 -818 3429
rect -784 3395 -778 3429
rect -824 3357 -778 3395
rect -824 3323 -818 3357
rect -784 3323 -778 3357
rect -824 3285 -778 3323
rect -824 3251 -818 3285
rect -784 3251 -778 3285
rect -824 3213 -778 3251
rect -824 3179 -818 3213
rect -784 3179 -778 3213
rect -824 3141 -778 3179
rect -68 3416 -62 3450
rect -28 3416 -22 3450
rect -68 3378 -22 3416
rect -68 3344 -62 3378
rect -28 3344 -22 3378
rect -68 3306 -22 3344
rect -68 3272 -62 3306
rect -28 3272 -22 3306
rect -68 3234 -22 3272
rect -68 3200 -62 3234
rect -28 3200 -22 3234
rect 161 3549 295 3561
rect 161 3515 167 3549
rect 201 3515 255 3549
rect 289 3515 295 3549
rect 161 3476 295 3515
rect 161 3442 167 3476
rect 201 3475 295 3476
rect 201 3442 255 3475
rect 161 3441 255 3442
rect 289 3441 295 3475
rect 161 3404 295 3441
rect 161 3370 167 3404
rect 201 3401 295 3404
rect 201 3370 255 3401
rect 161 3367 255 3370
rect 289 3367 295 3401
rect 161 3332 295 3367
rect 161 3298 167 3332
rect 201 3327 295 3332
rect 201 3298 255 3327
rect 161 3293 255 3298
rect 289 3293 295 3327
rect 161 3260 295 3293
rect 161 3226 167 3260
rect 201 3253 295 3260
rect 201 3226 255 3253
rect 161 3219 255 3226
rect 289 3219 295 3253
rect -68 3190 -22 3200
tri -22 3190 -4 3208 sw
rect -68 3160 -4 3190
tri -68 3154 -62 3160 ne
rect -62 3154 -4 3160
tri -62 3151 -59 3154 ne
rect -59 3151 -4 3154
tri -59 3142 -50 3151 ne
rect -824 3107 -818 3141
rect -784 3107 -778 3141
rect -824 3069 -778 3107
rect -824 3035 -818 3069
rect -784 3035 -778 3069
rect -824 2997 -778 3035
rect -824 2963 -818 2997
rect -784 2963 -778 2997
rect -824 2925 -778 2963
rect -824 2891 -818 2925
rect -784 2891 -778 2925
rect -824 2853 -778 2891
rect -824 2819 -818 2853
rect -784 2819 -778 2853
rect -824 2781 -778 2819
rect -824 2747 -818 2781
rect -784 2747 -778 2781
rect -824 2709 -778 2747
rect -824 2675 -818 2709
rect -784 2675 -778 2709
rect -824 2637 -778 2675
rect -824 2603 -818 2637
rect -784 2603 -778 2637
rect -824 2565 -778 2603
rect -824 2531 -818 2565
rect -784 2531 -778 2565
rect -824 2493 -778 2531
rect -824 2459 -818 2493
rect -784 2459 -778 2493
rect -824 2421 -778 2459
rect -824 2387 -818 2421
rect -784 2387 -778 2421
rect -824 2349 -778 2387
rect -824 2315 -818 2349
rect -784 2315 -778 2349
rect -824 2277 -778 2315
rect -824 2243 -818 2277
rect -784 2243 -778 2277
rect -824 2205 -778 2243
rect -824 2171 -818 2205
rect -784 2171 -778 2205
rect -824 2133 -778 2171
rect -824 2099 -818 2133
rect -784 2099 -778 2133
rect -824 2061 -778 2099
rect -824 2027 -818 2061
rect -784 2027 -778 2061
tri -830 2007 -824 2013 se
rect -824 2007 -778 2027
rect -830 2001 -778 2007
rect -830 1919 -778 1949
rect -830 1861 -778 1867
tri -830 1858 -827 1861 ne
rect -827 1858 -778 1861
tri -827 1857 -826 1858 ne
rect -826 1857 -778 1858
tri -826 1855 -824 1857 ne
rect -824 1845 -778 1857
rect -824 1811 -818 1845
rect -784 1811 -778 1845
rect -824 1773 -778 1811
rect -824 1739 -818 1773
rect -784 1739 -778 1773
rect -824 1701 -778 1739
rect -824 1667 -818 1701
rect -784 1667 -778 1701
rect -824 1629 -778 1667
rect -824 1595 -818 1629
rect -784 1595 -778 1629
rect -824 1557 -778 1595
rect -824 1523 -818 1557
rect -784 1523 -778 1557
rect -824 1485 -778 1523
rect -824 1451 -818 1485
rect -784 1451 -778 1485
rect -824 1413 -778 1451
rect -824 1379 -818 1413
rect -784 1379 -778 1413
rect -824 1341 -778 1379
rect -824 1307 -818 1341
rect -784 1307 -778 1341
rect -824 1269 -778 1307
rect -824 1235 -818 1269
rect -784 1235 -778 1269
rect -824 1197 -778 1235
rect -824 1163 -818 1197
rect -784 1163 -778 1197
rect -824 1125 -778 1163
rect -824 1091 -818 1125
rect -784 1091 -778 1125
rect -824 1053 -778 1091
rect -824 1019 -818 1053
rect -784 1019 -778 1053
rect -824 981 -778 1019
rect -824 947 -818 981
rect -784 947 -778 981
rect -824 909 -778 947
rect -824 875 -818 909
rect -784 875 -778 909
rect -824 837 -778 875
rect -824 803 -818 837
rect -784 803 -778 837
rect -824 765 -778 803
rect -824 731 -818 765
rect -784 731 -778 765
rect -824 693 -778 731
rect -824 659 -818 693
rect -784 659 -778 693
rect -824 621 -778 659
rect -824 587 -818 621
rect -784 587 -778 621
rect -824 548 -778 587
rect -824 514 -818 548
rect -784 514 -778 548
rect -824 475 -778 514
rect -824 441 -818 475
rect -784 441 -778 475
rect -824 402 -778 441
rect -824 368 -818 402
rect -784 368 -778 402
rect -824 329 -778 368
rect -824 295 -818 329
rect -784 295 -778 329
rect -824 256 -778 295
rect -824 222 -818 256
rect -784 222 -778 256
rect -824 183 -778 222
rect -824 149 -818 183
rect -784 149 -778 183
rect -824 110 -778 149
rect -824 76 -818 110
rect -784 76 -778 110
rect -824 37 -778 76
rect -824 3 -818 37
rect -784 3 -778 37
rect -824 -36 -778 3
rect -824 -70 -818 -36
rect -784 -70 -778 -36
rect -824 -109 -778 -70
rect -824 -143 -818 -109
rect -784 -143 -778 -109
rect -824 -182 -778 -143
rect -50 3117 -44 3151
rect -10 3117 -4 3151
rect -50 3079 -4 3117
rect -50 3045 -44 3079
rect -10 3045 -4 3079
rect -50 3007 -4 3045
rect -50 2973 -44 3007
rect -10 2973 -4 3007
rect -50 2935 -4 2973
rect -50 2901 -44 2935
rect -10 2901 -4 2935
rect -50 2863 -4 2901
rect -50 2829 -44 2863
rect -10 2829 -4 2863
rect -50 2791 -4 2829
rect -50 2757 -44 2791
rect -10 2757 -4 2791
rect -50 2719 -4 2757
rect -50 2685 -44 2719
rect -10 2685 -4 2719
rect -50 2647 -4 2685
rect -50 2613 -44 2647
rect -10 2613 -4 2647
rect -50 2575 -4 2613
rect -50 2541 -44 2575
rect -10 2541 -4 2575
rect -50 2503 -4 2541
rect -50 2469 -44 2503
rect -10 2469 -4 2503
rect -50 2431 -4 2469
rect -50 2397 -44 2431
rect -10 2397 -4 2431
rect -50 2359 -4 2397
rect -50 2325 -44 2359
rect -10 2325 -4 2359
rect -50 2287 -4 2325
rect -50 2253 -44 2287
rect -10 2253 -4 2287
rect -50 2215 -4 2253
rect -50 2181 -44 2215
rect -10 2181 -4 2215
rect -50 2143 -4 2181
rect -50 2109 -44 2143
rect -10 2109 -4 2143
rect -50 2071 -4 2109
rect -50 2037 -44 2071
rect -10 2037 -4 2071
rect -50 1999 -4 2037
rect -50 1965 -44 1999
rect -10 1965 -4 1999
rect -50 1927 -4 1965
rect -50 1893 -44 1927
rect -10 1893 -4 1927
rect -50 1855 -4 1893
rect -50 1821 -44 1855
rect -10 1821 -4 1855
rect -50 1783 -4 1821
rect -50 1749 -44 1783
rect -10 1749 -4 1783
rect -50 1711 -4 1749
rect -50 1677 -44 1711
rect -10 1677 -4 1711
rect -50 1639 -4 1677
rect -50 1605 -44 1639
rect -10 1605 -4 1639
rect -50 1567 -4 1605
rect -50 1533 -44 1567
rect -10 1533 -4 1567
rect -50 1495 -4 1533
rect -50 1461 -44 1495
rect -10 1461 -4 1495
rect -50 1423 -4 1461
rect -50 1389 -44 1423
rect -10 1389 -4 1423
rect -50 1351 -4 1389
rect -50 1317 -44 1351
rect -10 1317 -4 1351
rect -50 1279 -4 1317
rect -50 1245 -44 1279
rect -10 1245 -4 1279
rect -50 1207 -4 1245
rect -50 1173 -44 1207
rect -10 1173 -4 1207
rect -50 1135 -4 1173
rect -50 1101 -44 1135
rect -10 1101 -4 1135
rect -50 1063 -4 1101
rect -50 1029 -44 1063
rect -10 1029 -4 1063
rect -50 990 -4 1029
rect -50 956 -44 990
rect -10 956 -4 990
rect -50 917 -4 956
rect -50 883 -44 917
rect -10 883 -4 917
rect -50 844 -4 883
rect -50 810 -44 844
rect -10 810 -4 844
rect -50 771 -4 810
rect -50 737 -44 771
rect -10 737 -4 771
rect -50 698 -4 737
rect -50 664 -44 698
rect -10 664 -4 698
rect -50 625 -4 664
rect -50 591 -44 625
rect -10 591 -4 625
rect -50 552 -4 591
rect -50 518 -44 552
rect -10 518 -4 552
rect -50 479 -4 518
rect -50 445 -44 479
rect -10 445 -4 479
rect -50 406 -4 445
rect -50 372 -44 406
rect -10 372 -4 406
rect -50 333 -4 372
rect -50 299 -44 333
rect -10 299 -4 333
rect -50 260 -4 299
rect -50 226 -44 260
rect -10 236 -4 260
rect 161 3188 295 3219
rect 161 3154 167 3188
rect 201 3179 295 3188
rect 201 3154 255 3179
rect 161 3145 255 3154
rect 289 3145 295 3179
rect 161 3116 295 3145
rect 161 3082 167 3116
rect 201 3105 295 3116
rect 201 3082 255 3105
rect 161 3071 255 3082
rect 289 3071 295 3105
rect 161 3044 295 3071
rect 161 3010 167 3044
rect 201 3031 295 3044
rect 201 3010 255 3031
rect 161 2997 255 3010
rect 289 2997 295 3031
rect 161 2972 295 2997
rect 161 2938 167 2972
rect 201 2957 295 2972
rect 201 2938 255 2957
rect 161 2923 255 2938
rect 289 2923 295 2957
rect 161 2900 295 2923
rect 161 2866 167 2900
rect 201 2883 295 2900
rect 201 2866 255 2883
rect 161 2849 255 2866
rect 289 2849 295 2883
rect 161 2828 295 2849
rect 161 2794 167 2828
rect 201 2809 295 2828
rect 201 2794 255 2809
rect 161 2775 255 2794
rect 289 2775 295 2809
rect 161 2756 295 2775
rect 161 2722 167 2756
rect 201 2735 295 2756
rect 201 2722 255 2735
rect 161 2701 255 2722
rect 289 2701 295 2735
rect 161 2684 295 2701
rect 161 2650 167 2684
rect 201 2661 295 2684
rect 201 2650 255 2661
rect 161 2627 255 2650
rect 289 2627 295 2661
rect 161 2612 295 2627
rect 161 2578 167 2612
rect 201 2587 295 2612
rect 201 2578 255 2587
rect 161 2553 255 2578
rect 289 2553 295 2587
rect 161 2540 295 2553
rect 161 2506 167 2540
rect 201 2514 295 2540
rect 201 2506 255 2514
rect 161 2480 255 2506
rect 289 2480 295 2514
rect 161 2468 295 2480
rect 161 2434 167 2468
rect 201 2441 295 2468
rect 201 2434 255 2441
rect 161 2407 255 2434
rect 289 2407 295 2441
rect 161 2396 295 2407
rect 161 2362 167 2396
rect 201 2368 295 2396
rect 201 2362 255 2368
rect 161 2334 255 2362
rect 289 2334 295 2368
rect 161 2324 295 2334
rect 161 2290 167 2324
rect 201 2295 295 2324
rect 201 2290 255 2295
rect 161 2261 255 2290
rect 289 2261 295 2295
rect 161 2252 295 2261
rect 161 2218 167 2252
rect 201 2222 295 2252
rect 201 2218 255 2222
rect 161 2188 255 2218
rect 289 2188 295 2222
rect 161 2180 295 2188
rect 161 2146 167 2180
rect 201 2149 295 2180
rect 201 2146 255 2149
rect 161 2115 255 2146
rect 289 2115 295 2149
rect 161 2108 295 2115
rect 161 2074 167 2108
rect 201 2076 295 2108
rect 201 2074 255 2076
rect 161 2042 255 2074
rect 289 2042 295 2076
rect 161 2036 295 2042
rect 161 2002 167 2036
rect 201 2003 295 2036
rect 201 2002 255 2003
rect 161 1969 255 2002
rect 289 1969 295 2003
rect 161 1964 295 1969
rect 161 1930 167 1964
rect 201 1930 295 1964
rect 161 1896 255 1930
rect 289 1896 295 1930
rect 161 1892 295 1896
rect 161 1858 167 1892
rect 201 1858 295 1892
rect 161 1857 295 1858
rect 161 1823 255 1857
rect 289 1823 295 1857
rect 161 1820 295 1823
rect 161 1786 167 1820
rect 201 1786 295 1820
rect 161 1784 295 1786
rect 161 1750 255 1784
rect 289 1750 295 1784
rect 161 1748 295 1750
rect 161 1714 167 1748
rect 201 1714 295 1748
rect 161 1711 295 1714
rect 161 1677 255 1711
rect 289 1677 295 1711
rect 161 1676 295 1677
rect 161 1642 167 1676
rect 201 1642 295 1676
rect 161 1638 295 1642
rect 161 1604 255 1638
rect 289 1604 295 1638
rect 161 1570 167 1604
rect 201 1570 295 1604
rect 161 1565 295 1570
rect 161 1532 255 1565
rect 161 1498 167 1532
rect 201 1531 255 1532
rect 289 1531 295 1565
rect 201 1498 295 1531
rect 161 1492 295 1498
rect 161 1460 255 1492
rect 161 1426 167 1460
rect 201 1458 255 1460
rect 289 1458 295 1492
rect 201 1426 295 1458
rect 161 1419 295 1426
rect 161 1388 255 1419
rect 161 1354 167 1388
rect 201 1385 255 1388
rect 289 1385 295 1419
rect 201 1354 295 1385
rect 161 1346 295 1354
rect 161 1316 255 1346
rect 161 1282 167 1316
rect 201 1312 255 1316
rect 289 1312 295 1346
rect 201 1282 295 1312
rect 161 1273 295 1282
rect 161 1244 255 1273
rect 161 1210 167 1244
rect 201 1239 255 1244
rect 289 1239 295 1273
rect 201 1210 295 1239
rect 161 1200 295 1210
rect 161 1172 255 1200
rect 161 1138 167 1172
rect 201 1166 255 1172
rect 289 1166 295 1200
rect 201 1138 295 1166
rect 161 1127 295 1138
rect 161 1100 255 1127
rect 161 1066 167 1100
rect 201 1093 255 1100
rect 289 1093 295 1127
rect 201 1066 295 1093
rect 161 1054 295 1066
rect 161 1028 255 1054
rect 161 994 167 1028
rect 201 1020 255 1028
rect 289 1020 295 1054
rect 201 994 295 1020
rect 161 981 295 994
rect 161 956 255 981
rect 161 922 167 956
rect 201 947 255 956
rect 289 947 295 981
rect 201 922 295 947
rect 161 908 295 922
rect 161 884 255 908
rect 161 850 167 884
rect 201 874 255 884
rect 289 874 295 908
rect 201 850 295 874
rect 161 835 295 850
rect 161 812 255 835
rect 161 778 167 812
rect 201 801 255 812
rect 289 801 295 835
rect 201 778 295 801
rect 161 762 295 778
rect 161 740 255 762
rect 161 706 167 740
rect 201 728 255 740
rect 289 728 295 762
rect 201 706 295 728
rect 161 689 295 706
rect 161 668 255 689
rect 161 634 167 668
rect 201 655 255 668
rect 289 655 295 689
rect 201 634 295 655
rect 161 616 295 634
rect 161 596 255 616
rect 161 562 167 596
rect 201 582 255 596
rect 289 582 295 616
rect 201 562 295 582
rect 161 543 295 562
rect 161 524 255 543
rect 161 490 167 524
rect 201 509 255 524
rect 289 509 295 543
rect 201 490 295 509
rect 161 470 295 490
rect 161 452 255 470
rect 161 418 167 452
rect 201 436 255 452
rect 289 436 295 470
rect 364 3548 410 3587
rect 364 3514 370 3548
rect 404 3514 410 3548
rect 364 3475 410 3514
rect 364 3441 370 3475
rect 404 3441 410 3475
rect 364 3402 410 3441
rect 364 3368 370 3402
rect 404 3368 410 3402
rect 364 3329 410 3368
rect 364 3295 370 3329
rect 404 3295 410 3329
rect 364 3256 410 3295
rect 364 3222 370 3256
rect 404 3222 410 3256
rect 364 3183 410 3222
rect 364 3149 370 3183
rect 404 3149 410 3183
rect 364 3110 410 3149
rect 364 3076 370 3110
rect 404 3076 410 3110
rect 364 3037 410 3076
rect 364 3003 370 3037
rect 404 3003 410 3037
rect 364 2964 410 3003
rect 364 2930 370 2964
rect 404 2930 410 2964
rect 364 2891 410 2930
rect 364 2857 370 2891
rect 404 2857 410 2891
rect 364 2818 410 2857
rect 364 2784 370 2818
rect 404 2784 410 2818
rect 364 2745 410 2784
rect 364 2711 370 2745
rect 404 2711 410 2745
rect 364 2673 410 2711
rect 364 2639 370 2673
rect 404 2639 410 2673
rect 364 2601 410 2639
rect 364 2567 370 2601
rect 404 2567 410 2601
rect 364 2529 410 2567
rect 364 2495 370 2529
rect 404 2495 410 2529
rect 364 2457 410 2495
rect 364 2423 370 2457
rect 404 2423 410 2457
rect 364 2385 410 2423
rect 364 2351 370 2385
rect 404 2351 410 2385
rect 364 2313 410 2351
rect 364 2279 370 2313
rect 404 2279 410 2313
rect 364 2241 410 2279
rect 364 2207 370 2241
rect 404 2207 410 2241
rect 364 2169 410 2207
rect 364 2135 370 2169
rect 404 2135 410 2169
rect 364 2097 410 2135
rect 364 2063 370 2097
rect 404 2063 410 2097
rect 364 2016 410 2063
rect 364 1982 370 2016
rect 404 1982 410 2016
rect 364 1943 410 1982
rect 364 1909 370 1943
rect 404 1909 410 1943
rect 364 1870 410 1909
rect 364 1836 370 1870
rect 404 1836 410 1870
rect 364 1797 410 1836
rect 364 1763 370 1797
rect 404 1763 410 1797
rect 364 1725 410 1763
rect 364 1691 370 1725
rect 404 1691 410 1725
rect 364 1653 410 1691
rect 364 1619 370 1653
rect 404 1619 410 1653
rect 364 1581 410 1619
rect 364 1547 370 1581
rect 404 1547 410 1581
rect 364 1509 410 1547
rect 364 1475 370 1509
rect 404 1475 410 1509
rect 364 1437 410 1475
rect 364 1403 370 1437
rect 404 1403 410 1437
rect 364 1365 410 1403
rect 466 3659 512 3671
rect 466 3625 472 3659
rect 506 3625 512 3659
rect 466 3586 512 3625
rect 466 3552 472 3586
rect 506 3552 512 3586
rect 466 3513 512 3552
rect 466 3479 472 3513
rect 506 3479 512 3513
rect 466 3440 512 3479
rect 466 3406 472 3440
rect 506 3406 512 3440
rect 466 3367 512 3406
rect 466 3333 472 3367
rect 506 3333 512 3367
rect 466 3294 512 3333
rect 466 3260 472 3294
rect 506 3260 512 3294
rect 466 3221 512 3260
rect 466 3187 472 3221
rect 506 3187 512 3221
rect 466 3148 512 3187
rect 466 3114 472 3148
rect 506 3114 512 3148
rect 466 3074 512 3114
rect 466 3040 472 3074
rect 506 3040 512 3074
rect 466 3000 512 3040
rect 466 2966 472 3000
rect 506 2966 512 3000
rect 466 2926 512 2966
rect 466 2892 472 2926
rect 506 2892 512 2926
rect 466 2852 512 2892
rect 466 2818 472 2852
rect 506 2818 512 2852
rect 466 2778 512 2818
rect 466 2744 472 2778
rect 506 2744 512 2778
rect 466 2704 512 2744
rect 466 2670 472 2704
rect 506 2670 512 2704
rect 466 2630 512 2670
rect 466 2596 472 2630
rect 506 2596 512 2630
rect 466 2556 512 2596
rect 466 2522 472 2556
rect 506 2522 512 2556
rect 466 2482 512 2522
rect 466 2448 472 2482
rect 506 2448 512 2482
rect 466 2408 512 2448
rect 466 2374 472 2408
rect 506 2374 512 2408
rect 466 2334 512 2374
rect 466 2300 472 2334
rect 506 2300 512 2334
rect 466 2260 512 2300
rect 466 2226 472 2260
rect 506 2226 512 2260
rect 466 2186 512 2226
rect 466 2152 472 2186
rect 506 2152 512 2186
rect 466 2112 512 2152
rect 466 2078 472 2112
rect 506 2078 512 2112
rect 466 2038 512 2078
rect 466 2004 472 2038
rect 506 2004 512 2038
rect 466 1964 512 2004
rect 466 1930 472 1964
rect 506 1930 512 1964
rect 466 1890 512 1930
rect 633 3651 651 3685
rect 685 3651 703 3685
rect 633 3612 703 3651
rect 633 3578 651 3612
rect 685 3578 703 3612
rect 633 3539 703 3578
rect 633 3505 651 3539
rect 685 3505 703 3539
rect 633 3466 703 3505
rect 633 3432 651 3466
rect 685 3432 703 3466
rect 633 3393 703 3432
rect 633 3359 651 3393
rect 685 3359 703 3393
rect 633 3320 703 3359
rect 633 3286 651 3320
rect 685 3286 703 3320
rect 633 3247 703 3286
rect 633 3213 651 3247
rect 685 3213 703 3247
rect 633 3174 703 3213
rect 633 3140 651 3174
rect 685 3140 703 3174
rect 633 3101 703 3140
rect 633 3067 651 3101
rect 685 3067 703 3101
rect 633 3028 703 3067
rect 633 2994 651 3028
rect 685 2994 703 3028
rect 633 2955 703 2994
rect 633 2921 651 2955
rect 685 2921 703 2955
rect 633 2882 703 2921
rect 633 2848 651 2882
rect 685 2848 703 2882
rect 633 2809 703 2848
rect 633 2775 651 2809
rect 685 2775 703 2809
rect 633 2736 703 2775
rect 633 2702 651 2736
rect 685 2702 703 2736
rect 633 2663 703 2702
rect 633 2629 651 2663
rect 685 2629 703 2663
rect 633 2590 703 2629
rect 633 2556 651 2590
rect 685 2556 703 2590
rect 633 2517 703 2556
rect 633 2483 651 2517
rect 685 2483 703 2517
rect 633 2444 703 2483
rect 633 2410 651 2444
rect 685 2410 703 2444
rect 633 2371 703 2410
rect 633 2337 651 2371
rect 685 2337 703 2371
rect 633 2298 703 2337
rect 633 2264 651 2298
rect 685 2264 703 2298
rect 633 2225 703 2264
rect 633 2191 651 2225
rect 685 2191 703 2225
rect 633 2152 703 2191
rect 633 2118 651 2152
rect 685 2118 703 2152
rect 633 2079 703 2118
rect 633 2045 651 2079
rect 685 2045 703 2079
rect 633 2005 703 2045
tri 703 2005 796 2098 sw
rect 633 1924 796 2005
rect 633 1920 668 1924
tri 633 1891 662 1920 ne
rect 466 1856 472 1890
rect 506 1856 512 1890
rect 466 1816 512 1856
rect 466 1782 472 1816
rect 506 1782 512 1816
rect 466 1742 512 1782
rect 466 1708 472 1742
rect 506 1708 512 1742
rect 466 1668 512 1708
rect 466 1634 472 1668
rect 506 1634 512 1668
rect 466 1594 512 1634
rect 466 1560 472 1594
rect 506 1560 512 1594
rect 466 1520 512 1560
rect 466 1486 472 1520
rect 506 1486 512 1520
rect 466 1446 512 1486
rect 466 1412 472 1446
rect 506 1412 512 1446
rect 466 1400 512 1412
rect 662 1890 668 1920
rect 702 1890 756 1924
rect 790 1890 796 1924
rect 662 1852 796 1890
rect 662 1818 668 1852
rect 702 1851 796 1852
rect 702 1818 756 1851
rect 662 1817 756 1818
rect 790 1817 796 1851
rect 662 1780 796 1817
rect 662 1746 668 1780
rect 702 1778 796 1780
rect 702 1746 756 1778
rect 662 1744 756 1746
rect 790 1744 796 1778
rect 662 1708 796 1744
rect 662 1674 668 1708
rect 702 1705 796 1708
rect 702 1674 756 1705
rect 662 1671 756 1674
rect 790 1671 796 1705
rect 662 1636 796 1671
rect 662 1602 668 1636
rect 702 1632 796 1636
rect 702 1602 756 1632
rect 662 1598 756 1602
rect 790 1598 796 1632
rect 662 1564 796 1598
rect 662 1530 668 1564
rect 702 1559 796 1564
rect 702 1530 756 1559
rect 662 1525 756 1530
rect 790 1525 796 1559
rect 662 1492 796 1525
rect 662 1458 668 1492
rect 702 1486 796 1492
rect 702 1458 756 1486
rect 662 1452 756 1458
rect 790 1452 796 1486
rect 662 1419 796 1452
rect 886 1535 892 1587
rect 944 1535 961 1587
rect 1013 1535 1030 1587
rect 1082 1535 1088 1587
rect 886 1493 1088 1535
rect 886 1441 892 1493
rect 944 1441 961 1493
rect 1013 1441 1030 1493
rect 1082 1441 1088 1493
rect 364 1331 370 1365
rect 404 1331 410 1365
rect 364 1293 410 1331
rect 364 1259 370 1293
rect 404 1259 410 1293
rect 364 1221 410 1259
rect 364 1187 370 1221
rect 404 1187 410 1221
rect 364 1149 410 1187
rect 364 1115 370 1149
rect 404 1115 410 1149
rect 364 1077 410 1115
rect 364 1043 370 1077
rect 404 1043 410 1077
rect 364 1005 410 1043
rect 364 971 370 1005
rect 404 971 410 1005
rect 364 933 410 971
rect 364 899 370 933
rect 404 899 410 933
rect 364 861 410 899
rect 364 827 370 861
rect 404 827 410 861
rect 364 789 410 827
rect 364 755 370 789
rect 404 755 410 789
rect 364 717 410 755
rect 364 683 370 717
rect 404 683 410 717
rect 364 645 410 683
rect 364 611 370 645
rect 404 611 410 645
rect 364 573 410 611
rect 364 539 370 573
rect 404 539 410 573
rect 364 501 410 539
rect 364 467 370 501
rect 404 467 410 501
rect 364 455 410 467
rect 662 1385 668 1419
rect 702 1413 796 1419
rect 702 1385 756 1413
rect 662 1379 756 1385
rect 790 1379 796 1413
rect 662 1346 796 1379
rect 662 1312 668 1346
rect 702 1340 796 1346
rect 702 1312 756 1340
rect 662 1306 756 1312
rect 790 1306 796 1340
rect 662 1273 796 1306
rect 662 1239 668 1273
rect 702 1267 796 1273
rect 702 1239 756 1267
rect 662 1233 756 1239
rect 790 1233 796 1267
rect 662 1200 796 1233
rect 662 1166 668 1200
rect 702 1194 796 1200
rect 702 1166 756 1194
rect 662 1160 756 1166
rect 790 1160 796 1194
rect 662 1127 796 1160
rect 662 1093 668 1127
rect 702 1121 796 1127
rect 702 1093 756 1121
rect 662 1087 756 1093
rect 790 1087 796 1121
rect 662 1054 796 1087
rect 662 1020 668 1054
rect 702 1048 796 1054
rect 702 1020 756 1048
rect 662 1014 756 1020
rect 790 1014 796 1048
rect 662 981 796 1014
rect 662 947 668 981
rect 702 974 796 981
rect 702 947 756 974
rect 662 940 756 947
rect 790 940 796 974
rect 662 908 796 940
rect 662 874 668 908
rect 702 900 796 908
rect 702 874 756 900
rect 662 866 756 874
rect 790 866 796 900
rect 662 835 796 866
rect 662 801 668 835
rect 702 826 796 835
rect 702 801 756 826
rect 662 792 756 801
rect 790 792 796 826
rect 662 762 796 792
rect 662 728 668 762
rect 702 752 796 762
rect 702 728 756 752
rect 662 718 756 728
rect 790 718 796 752
rect 662 689 796 718
rect 662 655 668 689
rect 702 678 796 689
rect 702 655 756 678
rect 662 644 756 655
rect 790 644 796 678
rect 662 616 796 644
rect 662 582 668 616
rect 702 604 796 616
rect 702 582 756 604
rect 662 570 756 582
rect 790 570 796 604
rect 662 543 796 570
rect 662 509 668 543
rect 702 530 796 543
rect 702 509 756 530
rect 662 496 756 509
rect 790 496 796 530
rect 662 470 796 496
tri 295 436 296 437 sw
tri 661 436 662 437 se
rect 662 436 668 470
rect 702 456 796 470
rect 702 436 756 456
rect 201 422 296 436
tri 296 422 310 436 sw
tri 647 422 661 436 se
rect 661 422 756 436
rect 790 422 796 456
rect 201 418 310 422
rect 161 397 310 418
tri 310 397 335 422 sw
tri 622 397 647 422 se
rect 647 397 796 422
rect 161 380 255 397
rect 161 346 167 380
rect 201 363 255 380
rect 289 363 335 397
tri 335 363 369 397 sw
tri 588 363 622 397 se
rect 622 363 668 397
rect 702 382 796 397
rect 702 363 756 382
rect 201 348 369 363
tri 369 348 384 363 sw
tri 573 348 588 363 se
rect 588 348 756 363
rect 790 348 796 382
rect 201 346 384 348
rect 161 330 384 346
tri 384 330 402 348 sw
tri 555 330 573 348 se
rect 573 330 796 348
rect 161 324 796 330
rect 161 308 255 324
rect 161 274 167 308
rect 201 290 255 308
rect 289 290 338 324
rect 372 290 421 324
rect 455 290 504 324
rect 538 290 586 324
rect 620 290 668 324
rect 702 308 796 324
rect 702 290 756 308
rect 201 274 756 290
rect 790 274 796 308
tri -4 236 9 249 sw
rect 161 236 796 274
rect -10 226 9 236
rect -50 202 9 226
tri 9 202 43 236 sw
rect 161 202 239 236
rect 273 202 313 236
rect 347 202 387 236
rect 421 202 461 236
rect 495 202 535 236
rect 569 202 609 236
rect 643 202 683 236
rect 717 202 796 236
rect -50 196 43 202
tri 43 196 49 202 sw
rect 161 196 796 202
tri 836 196 886 246 se
rect -50 187 49 196
rect -50 153 -44 187
rect -10 153 49 187
rect -50 132 49 153
tri 49 132 113 196 sw
tri 772 132 836 196 se
rect 836 132 886 196
rect -50 114 113 132
rect -50 80 -44 114
rect -10 110 113 114
tri 113 110 135 132 sw
tri 750 110 772 132 se
rect 772 110 886 132
tri 886 110 908 132 se
rect 908 110 936 132
rect -10 103 135 110
tri 135 103 142 110 sw
tri 743 103 750 110 se
rect 750 103 936 110
rect -10 95 936 103
rect -10 80 59 95
rect -50 61 59 80
rect 93 61 134 95
rect 168 61 209 95
rect 243 61 284 95
rect 318 61 359 95
rect 393 61 434 95
rect 468 61 509 95
rect 543 61 584 95
rect 618 61 659 95
rect 693 61 734 95
rect 768 61 808 95
rect 842 61 936 95
rect -50 41 936 61
rect -50 7 -44 41
rect -10 19 936 41
rect -10 7 36 19
rect -50 -15 36 7
rect 70 -15 113 19
rect 147 -15 190 19
rect 224 -15 267 19
rect 301 -15 344 19
rect 378 -15 421 19
rect 455 -15 498 19
rect 532 -15 575 19
rect 609 -15 653 19
rect 687 -15 731 19
rect 765 -15 809 19
rect 843 -15 936 19
rect -50 -54 936 -15
rect -50 -65 886 -54
rect -50 -99 36 -65
rect 70 -99 113 -65
rect 147 -99 190 -65
rect 224 -99 267 -65
rect 301 -99 344 -65
rect 378 -99 421 -65
rect 455 -99 498 -65
rect 532 -99 575 -65
rect 609 -99 653 -65
rect 687 -99 731 -65
rect 765 -99 809 -65
rect 843 -99 886 -65
tri 886 -76 908 -54 ne
rect 908 -76 936 -54
rect -50 -149 886 -99
rect -824 -216 -818 -182
rect -784 -183 -778 -182
tri -778 -183 -748 -153 sw
rect -50 -183 36 -149
rect 70 -183 113 -149
rect 147 -183 190 -149
rect 224 -183 267 -149
rect 301 -183 344 -149
rect 378 -183 421 -149
rect 455 -183 498 -149
rect 532 -183 575 -149
rect 609 -183 653 -149
rect 687 -183 731 -149
rect 765 -183 809 -149
rect 843 -183 886 -149
rect -784 -203 -748 -183
tri -748 -203 -728 -183 sw
rect -784 -215 -728 -203
tri -728 -215 -716 -203 sw
rect -50 -215 886 -183
rect -784 -216 -716 -215
rect -824 -243 -716 -216
tri -716 -243 -688 -215 sw
rect -824 -249 -688 -243
tri -688 -249 -682 -243 sw
rect -50 -249 -42 -215
rect -8 -233 886 -215
rect -8 -249 36 -233
rect -824 -255 -682 -249
rect -824 -289 -818 -255
rect -784 -289 -730 -255
rect -696 -267 -682 -255
tri -682 -267 -664 -249 sw
rect -50 -267 36 -249
rect 70 -267 113 -233
rect 147 -267 190 -233
rect 224 -267 267 -233
rect 301 -267 344 -233
rect 378 -267 421 -233
rect 455 -267 498 -233
rect 532 -267 575 -233
rect 609 -267 653 -233
rect 687 -267 731 -233
rect 765 -267 809 -233
rect 843 -267 886 -233
rect -696 -281 -664 -267
tri -664 -281 -650 -267 sw
rect -50 -281 886 -267
rect -696 -287 -650 -281
tri -650 -287 -644 -281 sw
rect -126 -287 886 -281
rect -696 -289 -644 -287
rect -824 -321 -644 -289
tri -644 -321 -610 -287 sw
rect -126 -321 -114 -287
rect -80 -321 -42 -287
rect -8 -317 886 -287
rect -8 -321 36 -317
rect -824 -327 -610 -321
tri -610 -327 -604 -321 sw
rect -126 -327 36 -321
rect -824 -361 -730 -327
rect -696 -333 -604 -327
tri -604 -333 -598 -327 sw
rect -696 -351 -598 -333
tri -598 -351 -580 -333 sw
rect -50 -351 36 -327
rect 70 -351 113 -317
rect 147 -351 190 -317
rect 224 -351 267 -317
rect 301 -351 344 -317
rect 378 -351 421 -317
rect 455 -351 498 -317
rect 532 -351 575 -317
rect 609 -351 653 -317
rect 687 -351 731 -317
rect 765 -351 809 -317
rect 843 -351 886 -317
rect -696 -361 -580 -351
rect -824 -363 -580 -361
tri -580 -363 -568 -351 sw
rect -824 -376 -803 -363
rect -736 -373 -690 -363
rect -50 -364 886 -351
tri -824 -397 -803 -376 ne
<< via1 >>
rect -830 14013 -778 14029
rect -830 13979 -818 14013
rect -818 13979 -784 14013
rect -784 13979 -778 14013
rect -830 13977 -778 13979
rect -830 13941 -778 13955
rect -830 13907 -818 13941
rect -818 13907 -784 13941
rect -784 13907 -778 13941
rect -830 13903 -778 13907
rect -830 13869 -778 13881
rect -830 13835 -818 13869
rect -818 13835 -784 13869
rect -784 13835 -778 13869
rect -830 13829 -778 13835
rect -830 13797 -778 13807
rect -830 13763 -818 13797
rect -818 13763 -784 13797
rect -784 13763 -778 13797
rect -830 13755 -778 13763
rect -830 13725 -778 13733
rect -830 13691 -818 13725
rect -818 13691 -784 13725
rect -784 13691 -778 13725
rect -830 13681 -778 13691
rect -310 14001 -258 14027
rect -310 13975 -305 14001
rect -305 13975 -271 14001
rect -271 13975 -258 14001
rect -242 14001 -190 14027
rect -242 13975 -231 14001
rect -231 13975 -197 14001
rect -197 13975 -190 14001
rect -174 14001 -122 14027
rect -174 13975 -157 14001
rect -157 13975 -123 14001
rect -123 13975 -122 14001
rect -310 13929 -258 13930
rect -310 13895 -305 13929
rect -305 13895 -271 13929
rect -271 13895 -258 13929
rect -310 13878 -258 13895
rect -242 13929 -190 13930
rect -242 13895 -231 13929
rect -231 13895 -197 13929
rect -197 13895 -190 13929
rect -242 13878 -190 13895
rect -174 13929 -122 13930
rect -174 13895 -157 13929
rect -157 13895 -123 13929
rect -123 13895 -122 13929
rect -174 13878 -122 13895
rect -310 13823 -305 13833
rect -305 13823 -271 13833
rect -271 13823 -258 13833
rect -310 13785 -258 13823
rect -310 13781 -305 13785
rect -305 13781 -271 13785
rect -271 13781 -258 13785
rect -242 13823 -231 13833
rect -231 13823 -197 13833
rect -197 13823 -190 13833
rect -242 13785 -190 13823
rect -242 13781 -231 13785
rect -231 13781 -197 13785
rect -197 13781 -190 13785
rect -174 13823 -157 13833
rect -157 13823 -123 13833
rect -123 13823 -122 13833
rect -174 13785 -122 13823
rect -174 13781 -157 13785
rect -157 13781 -123 13785
rect -123 13781 -122 13785
rect -310 13713 -258 13735
rect -310 13683 -305 13713
rect -305 13683 -271 13713
rect -271 13683 -258 13713
rect -242 13713 -190 13735
rect -242 13683 -231 13713
rect -231 13683 -197 13713
rect -197 13683 -190 13713
rect -174 13713 -122 13735
rect -174 13683 -157 13713
rect -157 13683 -123 13713
rect -123 13683 -122 13713
rect 216 14024 268 14029
rect 216 13990 245 14024
rect 245 13990 268 14024
rect 216 13977 268 13990
rect 281 14024 333 14029
rect 281 13990 293 14024
rect 293 13990 327 14024
rect 327 13990 333 14024
rect 281 13977 333 13990
rect 347 14024 399 14029
rect 413 14024 465 14029
rect 479 14024 531 14029
rect 545 14024 597 14029
rect 347 13990 375 14024
rect 375 13990 399 14024
rect 413 13990 457 14024
rect 457 13990 465 14024
rect 479 13990 491 14024
rect 491 13990 531 14024
rect 545 13990 573 14024
rect 573 13990 597 14024
rect 347 13977 399 13990
rect 413 13977 465 13990
rect 479 13977 531 13990
rect 545 13977 597 13990
rect 611 14024 663 14029
rect 611 13990 621 14024
rect 621 13990 655 14024
rect 655 13990 663 14024
rect 611 13977 663 13990
rect 677 14024 729 14029
rect 677 13990 703 14024
rect 703 13990 729 14024
rect 677 13977 729 13990
rect 216 13951 268 13955
rect 216 13917 245 13951
rect 245 13917 268 13951
rect 216 13903 268 13917
rect 281 13951 333 13955
rect 281 13917 293 13951
rect 293 13917 327 13951
rect 327 13917 333 13951
rect 281 13903 333 13917
rect 347 13951 399 13955
rect 413 13951 465 13955
rect 479 13951 531 13955
rect 545 13951 597 13955
rect 347 13917 375 13951
rect 375 13917 399 13951
rect 413 13917 457 13951
rect 457 13917 465 13951
rect 479 13917 491 13951
rect 491 13917 531 13951
rect 545 13917 573 13951
rect 573 13917 597 13951
rect 347 13903 399 13917
rect 413 13903 465 13917
rect 479 13903 531 13917
rect 545 13903 597 13917
rect 611 13951 663 13955
rect 611 13917 621 13951
rect 621 13917 655 13951
rect 655 13917 663 13951
rect 611 13903 663 13917
rect 677 13951 729 13955
rect 677 13917 703 13951
rect 703 13917 729 13951
rect 677 13903 729 13917
rect 216 13878 268 13881
rect 216 13844 245 13878
rect 245 13844 268 13878
rect 216 13829 268 13844
rect 281 13878 333 13881
rect 281 13844 293 13878
rect 293 13844 327 13878
rect 327 13844 333 13878
rect 281 13829 333 13844
rect 347 13878 399 13881
rect 413 13878 465 13881
rect 479 13878 531 13881
rect 545 13878 597 13881
rect 347 13844 375 13878
rect 375 13844 399 13878
rect 413 13844 457 13878
rect 457 13844 465 13878
rect 479 13844 491 13878
rect 491 13844 531 13878
rect 545 13844 573 13878
rect 573 13844 597 13878
rect 347 13829 399 13844
rect 413 13829 465 13844
rect 479 13829 531 13844
rect 545 13829 597 13844
rect 611 13878 663 13881
rect 611 13844 621 13878
rect 621 13844 655 13878
rect 655 13844 663 13878
rect 611 13829 663 13844
rect 677 13878 729 13881
rect 677 13844 703 13878
rect 703 13844 729 13878
rect 677 13829 729 13844
rect 216 13805 268 13807
rect 216 13771 245 13805
rect 245 13771 268 13805
rect 216 13755 268 13771
rect 281 13805 333 13807
rect 281 13771 293 13805
rect 293 13771 327 13805
rect 327 13771 333 13805
rect 281 13755 333 13771
rect 347 13805 399 13807
rect 413 13805 465 13807
rect 479 13805 531 13807
rect 545 13805 597 13807
rect 347 13771 375 13805
rect 375 13771 399 13805
rect 413 13771 457 13805
rect 457 13771 465 13805
rect 479 13771 491 13805
rect 491 13771 531 13805
rect 545 13771 573 13805
rect 573 13771 597 13805
rect 347 13755 399 13771
rect 413 13755 465 13771
rect 479 13755 531 13771
rect 545 13755 597 13771
rect 611 13805 663 13807
rect 611 13771 621 13805
rect 621 13771 655 13805
rect 655 13771 663 13805
rect 611 13755 663 13771
rect 677 13805 729 13807
rect 677 13771 703 13805
rect 703 13771 729 13805
rect 677 13755 729 13771
rect 216 13732 268 13733
rect 216 13698 245 13732
rect 245 13698 268 13732
rect 216 13681 268 13698
rect 281 13732 333 13733
rect 281 13698 293 13732
rect 293 13698 327 13732
rect 327 13698 333 13732
rect 281 13681 333 13698
rect 347 13732 399 13733
rect 413 13732 465 13733
rect 479 13732 531 13733
rect 545 13732 597 13733
rect 347 13698 375 13732
rect 375 13698 399 13732
rect 413 13698 457 13732
rect 457 13698 465 13732
rect 479 13698 491 13732
rect 491 13698 531 13732
rect 545 13698 573 13732
rect 573 13698 597 13732
rect 347 13681 399 13698
rect 413 13681 465 13698
rect 479 13681 531 13698
rect 545 13681 597 13698
rect 611 13732 663 13733
rect 611 13698 621 13732
rect 621 13698 655 13732
rect 655 13698 663 13732
rect 611 13681 663 13698
rect 677 13732 729 13733
rect 677 13698 703 13732
rect 703 13698 729 13732
rect 677 13681 729 13698
rect 887 13977 939 14029
rect 961 13977 1013 14029
rect 1035 13977 1087 14029
rect 887 13903 939 13955
rect 961 13903 1013 13955
rect 1035 13903 1087 13955
rect 887 13829 939 13881
rect 961 13829 1013 13881
rect 1035 13829 1087 13881
rect 887 13755 939 13807
rect 961 13755 1013 13807
rect 1035 13755 1087 13807
rect 887 13681 939 13733
rect 961 13681 1013 13733
rect 1035 13681 1087 13733
rect -305 12129 -253 12166
rect -305 12114 -271 12129
rect -271 12114 -253 12129
rect -240 12129 -188 12166
rect -240 12114 -231 12129
rect -231 12114 -197 12129
rect -197 12114 -188 12129
rect -175 12129 -123 12166
rect -175 12114 -157 12129
rect -157 12114 -123 12129
rect -62 12114 -10 12166
rect 8 12114 60 12166
rect 78 12114 130 12166
rect 148 12114 200 12166
rect 218 12114 270 12166
rect 289 12114 341 12166
rect -310 6382 -305 6391
rect -305 6382 -271 6391
rect -271 6382 -258 6391
rect -310 6343 -258 6382
rect -310 6339 -305 6343
rect -305 6339 -271 6343
rect -271 6339 -258 6343
rect -240 6382 -231 6391
rect -231 6382 -197 6391
rect -197 6382 -188 6391
rect -240 6343 -188 6382
rect -240 6339 -231 6343
rect -231 6339 -197 6343
rect -197 6339 -188 6343
rect -170 6382 -157 6391
rect -157 6382 -123 6391
rect -123 6382 -118 6391
rect -170 6343 -118 6382
rect -170 6339 -157 6343
rect -157 6339 -123 6343
rect -123 6339 -118 6343
rect -310 6309 -305 6321
rect -305 6309 -271 6321
rect -271 6309 -258 6321
rect -310 6270 -258 6309
rect -310 6269 -305 6270
rect -305 6269 -271 6270
rect -271 6269 -258 6270
rect -240 6309 -231 6321
rect -231 6309 -197 6321
rect -197 6309 -188 6321
rect -240 6270 -188 6309
rect -240 6269 -231 6270
rect -231 6269 -197 6270
rect -197 6269 -188 6270
rect -170 6309 -157 6321
rect -157 6309 -123 6321
rect -123 6309 -118 6321
rect -170 6270 -118 6309
rect -170 6269 -157 6270
rect -157 6269 -123 6270
rect -123 6269 -118 6270
rect -310 6236 -305 6251
rect -305 6236 -271 6251
rect -271 6236 -258 6251
rect -310 6199 -258 6236
rect -240 6236 -231 6251
rect -231 6236 -197 6251
rect -197 6236 -188 6251
rect -240 6199 -188 6236
rect -170 6236 -157 6251
rect -157 6236 -123 6251
rect -123 6236 -118 6251
rect -170 6199 -118 6236
rect -310 6163 -305 6181
rect -305 6163 -271 6181
rect -271 6163 -258 6181
rect -310 6129 -258 6163
rect -240 6163 -231 6181
rect -231 6163 -197 6181
rect -197 6163 -188 6181
rect -240 6129 -188 6163
rect -170 6163 -157 6181
rect -157 6163 -123 6181
rect -123 6163 -118 6181
rect -170 6129 -118 6163
rect -310 6090 -305 6111
rect -305 6090 -271 6111
rect -271 6090 -258 6111
rect -310 6059 -258 6090
rect -240 6090 -231 6111
rect -231 6090 -197 6111
rect -197 6090 -188 6111
rect -240 6059 -188 6090
rect -170 6090 -157 6111
rect -157 6090 -123 6111
rect -123 6090 -118 6111
rect -170 6059 -118 6090
rect -310 6017 -305 6041
rect -305 6017 -271 6041
rect -271 6017 -258 6041
rect -310 5989 -258 6017
rect -240 6017 -231 6041
rect -231 6017 -197 6041
rect -197 6017 -188 6041
rect -240 5989 -188 6017
rect -170 6017 -157 6041
rect -157 6017 -123 6041
rect -123 6017 -118 6041
rect -170 5989 -118 6017
rect -310 5944 -305 5971
rect -305 5944 -271 5971
rect -271 5944 -258 5971
rect -310 5919 -258 5944
rect -240 5944 -231 5971
rect -231 5944 -197 5971
rect -197 5944 -188 5971
rect -240 5919 -188 5944
rect -170 5944 -157 5971
rect -157 5944 -123 5971
rect -123 5944 -118 5971
rect -170 5919 -118 5944
rect -310 5871 -305 5901
rect -305 5871 -271 5901
rect -271 5871 -258 5901
rect -310 5849 -258 5871
rect -240 5871 -231 5901
rect -231 5871 -197 5901
rect -197 5871 -188 5901
rect -240 5849 -188 5871
rect -170 5871 -157 5901
rect -157 5871 -123 5901
rect -123 5871 -118 5901
rect -170 5849 -118 5871
rect -310 5798 -305 5830
rect -305 5798 -271 5830
rect -271 5798 -258 5830
rect -310 5778 -258 5798
rect -240 5798 -231 5830
rect -231 5798 -197 5830
rect -197 5798 -188 5830
rect -240 5778 -188 5798
rect -170 5798 -157 5830
rect -157 5798 -123 5830
rect -123 5798 -118 5830
rect -170 5778 -118 5798
rect -68 6339 -16 6391
rect -68 6269 -16 6321
rect -68 6199 -16 6251
rect -68 6129 -16 6181
rect -68 6059 -16 6111
rect -68 5989 -16 6041
rect -68 5919 -16 5971
rect -68 5849 -16 5901
rect -68 5778 -16 5830
rect -310 5068 -305 5070
rect -305 5068 -271 5070
rect -271 5068 -258 5070
rect -310 5029 -258 5068
rect -310 5018 -305 5029
rect -305 5018 -271 5029
rect -271 5018 -258 5029
rect -240 5068 -231 5070
rect -231 5068 -197 5070
rect -197 5068 -188 5070
rect -240 5029 -188 5068
rect -240 5018 -231 5029
rect -231 5018 -197 5029
rect -197 5018 -188 5029
rect -170 5068 -157 5070
rect -157 5068 -123 5070
rect -123 5068 -118 5070
rect -170 5029 -118 5068
rect -170 5018 -157 5029
rect -157 5018 -123 5029
rect -123 5018 -118 5029
rect -310 4995 -305 5004
rect -305 4995 -271 5004
rect -271 4995 -258 5004
rect -310 4956 -258 4995
rect -310 4952 -305 4956
rect -305 4952 -271 4956
rect -271 4952 -258 4956
rect -240 4995 -231 5004
rect -231 4995 -197 5004
rect -197 4995 -188 5004
rect -240 4956 -188 4995
rect -240 4952 -231 4956
rect -231 4952 -197 4956
rect -197 4952 -188 4956
rect -170 4995 -157 5004
rect -157 4995 -123 5004
rect -123 4995 -118 5004
rect -170 4956 -118 4995
rect -170 4952 -157 4956
rect -157 4952 -123 4956
rect -123 4952 -118 4956
rect -310 4922 -305 4938
rect -305 4922 -271 4938
rect -271 4922 -258 4938
rect -310 4886 -258 4922
rect -240 4922 -231 4938
rect -231 4922 -197 4938
rect -197 4922 -188 4938
rect -240 4886 -188 4922
rect -170 4922 -157 4938
rect -157 4922 -123 4938
rect -123 4922 -118 4938
rect -170 4886 -118 4922
rect -310 4849 -305 4872
rect -305 4849 -271 4872
rect -271 4849 -258 4872
rect -310 4820 -258 4849
rect -240 4849 -231 4872
rect -231 4849 -197 4872
rect -197 4849 -188 4872
rect -240 4820 -188 4849
rect -170 4849 -157 4872
rect -157 4849 -123 4872
rect -123 4849 -118 4872
rect -170 4820 -118 4849
rect -310 4776 -305 4806
rect -305 4776 -271 4806
rect -271 4776 -258 4806
rect -310 4754 -258 4776
rect -240 4776 -231 4806
rect -231 4776 -197 4806
rect -197 4776 -188 4806
rect -240 4754 -188 4776
rect -170 4776 -157 4806
rect -157 4776 -123 4806
rect -123 4776 -118 4806
rect -170 4754 -118 4776
rect -310 4737 -258 4740
rect -310 4703 -305 4737
rect -305 4703 -271 4737
rect -271 4703 -258 4737
rect -310 4688 -258 4703
rect -240 4737 -188 4740
rect -240 4703 -231 4737
rect -231 4703 -197 4737
rect -197 4703 -188 4737
rect -240 4688 -188 4703
rect -170 4737 -118 4740
rect -170 4703 -157 4737
rect -157 4703 -123 4737
rect -123 4703 -118 4737
rect -170 4688 -118 4703
rect -310 4664 -258 4674
rect -310 4630 -305 4664
rect -305 4630 -271 4664
rect -271 4630 -258 4664
rect -310 4622 -258 4630
rect -240 4664 -188 4674
rect -240 4630 -231 4664
rect -231 4630 -197 4664
rect -197 4630 -188 4664
rect -240 4622 -188 4630
rect -170 4664 -118 4674
rect -170 4630 -157 4664
rect -157 4630 -123 4664
rect -123 4630 -118 4664
rect -170 4622 -118 4630
rect -310 4591 -258 4607
rect -310 4557 -305 4591
rect -305 4557 -271 4591
rect -271 4557 -258 4591
rect -310 4555 -258 4557
rect -240 4591 -188 4607
rect -240 4557 -231 4591
rect -231 4557 -197 4591
rect -197 4557 -188 4591
rect -240 4555 -188 4557
rect -170 4591 -118 4607
rect -170 4557 -157 4591
rect -157 4557 -123 4591
rect -123 4557 -118 4591
rect -170 4555 -118 4557
rect -310 4518 -258 4540
rect -310 4488 -305 4518
rect -305 4488 -271 4518
rect -271 4488 -258 4518
rect -240 4518 -188 4540
rect -240 4488 -231 4518
rect -231 4488 -197 4518
rect -197 4488 -188 4518
rect -170 4518 -118 4540
rect -170 4488 -157 4518
rect -157 4488 -123 4518
rect -123 4488 -118 4518
rect -310 4445 -258 4473
rect -310 4421 -305 4445
rect -305 4421 -271 4445
rect -271 4421 -258 4445
rect -240 4445 -188 4473
rect -240 4421 -231 4445
rect -231 4421 -197 4445
rect -197 4421 -188 4445
rect -170 4445 -118 4473
rect -170 4421 -157 4445
rect -157 4421 -123 4445
rect -123 4421 -118 4445
rect -310 4372 -258 4406
rect -310 4354 -305 4372
rect -305 4354 -271 4372
rect -271 4354 -258 4372
rect -240 4372 -188 4406
rect -240 4354 -231 4372
rect -231 4354 -197 4372
rect -197 4354 -188 4372
rect -170 4372 -118 4406
rect -170 4354 -157 4372
rect -157 4354 -123 4372
rect -123 4354 -118 4372
rect -310 4338 -305 4339
rect -305 4338 -271 4339
rect -271 4338 -258 4339
rect -310 4299 -258 4338
rect -310 4287 -305 4299
rect -305 4287 -271 4299
rect -271 4287 -258 4299
rect -240 4338 -231 4339
rect -231 4338 -197 4339
rect -197 4338 -188 4339
rect -240 4299 -188 4338
rect -240 4287 -231 4299
rect -231 4287 -197 4299
rect -197 4287 -188 4299
rect -170 4338 -157 4339
rect -157 4338 -123 4339
rect -123 4338 -118 4339
rect -170 4299 -118 4338
rect -170 4287 -157 4299
rect -157 4287 -123 4299
rect -123 4287 -118 4299
rect -310 4265 -305 4272
rect -305 4265 -271 4272
rect -271 4265 -258 4272
rect -310 4226 -258 4265
rect -310 4220 -305 4226
rect -305 4220 -271 4226
rect -271 4220 -258 4226
rect -240 4265 -231 4272
rect -231 4265 -197 4272
rect -197 4265 -188 4272
rect -240 4226 -188 4265
rect -240 4220 -231 4226
rect -231 4220 -197 4226
rect -197 4220 -188 4226
rect -170 4265 -157 4272
rect -157 4265 -123 4272
rect -123 4265 -118 4272
rect -170 4226 -118 4265
rect -170 4220 -157 4226
rect -157 4220 -123 4226
rect -123 4220 -118 4226
rect -310 4192 -305 4205
rect -305 4192 -271 4205
rect -271 4192 -258 4205
rect -310 4153 -258 4192
rect -240 4192 -231 4205
rect -231 4192 -197 4205
rect -197 4192 -188 4205
rect -240 4153 -188 4192
rect -170 4192 -157 4205
rect -157 4192 -123 4205
rect -123 4192 -118 4205
rect -170 4153 -118 4192
rect -310 4119 -305 4138
rect -305 4119 -271 4138
rect -271 4119 -258 4138
rect -310 4086 -258 4119
rect -240 4119 -231 4138
rect -231 4119 -197 4138
rect -197 4119 -188 4138
rect -240 4086 -188 4119
rect -170 4119 -157 4138
rect -157 4119 -123 4138
rect -123 4119 -118 4138
rect -170 4086 -118 4119
rect -310 4046 -305 4071
rect -305 4046 -271 4071
rect -271 4046 -258 4071
rect -310 4019 -258 4046
rect -240 4046 -231 4071
rect -231 4046 -197 4071
rect -197 4046 -188 4071
rect -240 4019 -188 4046
rect -170 4046 -157 4071
rect -157 4046 -123 4071
rect -123 4046 -118 4071
rect -170 4019 -118 4046
rect -68 5018 -16 5070
rect -68 4974 -16 5004
rect -68 4952 -62 4974
rect -62 4952 -28 4974
rect -28 4952 -16 4974
rect -68 4901 -16 4938
rect -68 4886 -62 4901
rect -62 4886 -28 4901
rect -28 4886 -16 4901
rect -68 4867 -62 4872
rect -62 4867 -28 4872
rect -28 4867 -16 4872
rect -68 4828 -16 4867
rect -68 4820 -62 4828
rect -62 4820 -28 4828
rect -28 4820 -16 4828
rect -68 4794 -62 4806
rect -62 4794 -28 4806
rect -28 4794 -16 4806
rect -68 4755 -16 4794
rect -68 4754 -62 4755
rect -62 4754 -28 4755
rect -28 4754 -16 4755
rect -68 4721 -62 4740
rect -62 4721 -28 4740
rect -28 4721 -16 4740
rect -68 4688 -16 4721
rect -68 4648 -62 4674
rect -62 4648 -28 4674
rect -28 4648 -16 4674
rect -68 4622 -16 4648
rect -68 4575 -62 4607
rect -62 4575 -28 4607
rect -28 4575 -16 4607
rect -68 4555 -16 4575
rect -68 4536 -16 4540
rect -68 4502 -62 4536
rect -62 4502 -28 4536
rect -28 4502 -16 4536
rect -68 4488 -16 4502
rect -68 4463 -16 4473
rect -68 4429 -62 4463
rect -62 4429 -28 4463
rect -28 4429 -16 4463
rect -68 4421 -16 4429
rect -68 4390 -16 4406
rect -68 4356 -62 4390
rect -62 4356 -28 4390
rect -28 4356 -16 4390
rect -68 4354 -16 4356
rect -68 4317 -16 4339
rect -68 4287 -62 4317
rect -62 4287 -28 4317
rect -28 4287 -16 4317
rect -68 4244 -16 4272
rect -68 4220 -62 4244
rect -62 4220 -28 4244
rect -28 4220 -16 4244
rect -68 4171 -16 4205
rect -68 4153 -62 4171
rect -62 4153 -28 4171
rect -28 4153 -16 4171
rect -68 4137 -62 4138
rect -62 4137 -28 4138
rect -28 4137 -16 4138
rect -68 4098 -16 4137
rect -68 4086 -62 4098
rect -62 4086 -28 4098
rect -28 4086 -16 4098
rect -68 4064 -62 4071
rect -62 4064 -28 4071
rect -28 4064 -16 4071
rect -68 4026 -16 4064
rect -68 4019 -62 4026
rect -62 4019 -28 4026
rect -28 4019 -16 4026
rect 162 4668 171 4691
rect 171 4668 205 4691
rect 205 4668 214 4691
rect 162 4639 214 4668
rect 162 4592 171 4625
rect 171 4592 205 4625
rect 205 4592 214 4625
rect 162 4573 214 4592
rect 162 4550 214 4558
rect 162 4516 171 4550
rect 171 4516 205 4550
rect 205 4516 214 4550
rect 162 4506 214 4516
rect 162 4474 214 4491
rect 162 4440 171 4474
rect 171 4440 205 4474
rect 205 4440 214 4474
rect 162 4439 214 4440
rect 162 4398 214 4424
rect 162 4372 171 4398
rect 171 4372 205 4398
rect 205 4372 214 4398
rect 162 4322 214 4357
rect 162 4305 171 4322
rect 171 4305 205 4322
rect 205 4305 214 4322
rect 162 4288 171 4290
rect 171 4288 205 4290
rect 205 4288 214 4290
rect 162 4246 214 4288
rect 162 4238 171 4246
rect 171 4238 205 4246
rect 205 4238 214 4246
rect 162 4212 171 4223
rect 171 4212 205 4223
rect 205 4212 214 4223
rect 162 4171 214 4212
rect -830 1989 -778 2001
rect -830 1955 -818 1989
rect -818 1955 -784 1989
rect -784 1955 -778 1989
rect -830 1949 -778 1955
rect -830 1917 -778 1919
rect -830 1883 -818 1917
rect -818 1883 -784 1917
rect -784 1883 -778 1917
rect -830 1867 -778 1883
rect 892 1535 944 1587
rect 961 1535 1013 1587
rect 1030 1535 1082 1587
rect 892 1441 944 1493
rect 961 1441 1013 1493
rect 1030 1441 1082 1493
<< metal2 >>
rect -830 14029 1088 14035
rect -778 14027 216 14029
rect -778 13977 -310 14027
rect -830 13975 -310 13977
rect -258 13975 -242 14027
rect -190 13975 -174 14027
rect -122 13977 216 14027
rect 268 13977 281 14029
rect 333 13977 347 14029
rect 399 13977 413 14029
rect 465 13977 479 14029
rect 531 13977 545 14029
rect 597 13977 611 14029
rect 663 13977 677 14029
rect 729 13977 887 14029
rect 939 13977 961 14029
rect 1013 13977 1035 14029
rect 1087 13977 1088 14029
rect -122 13975 1088 13977
rect -830 13955 1088 13975
rect -778 13930 216 13955
rect -778 13903 -310 13930
rect -830 13881 -310 13903
rect -778 13878 -310 13881
rect -258 13878 -242 13930
rect -190 13878 -174 13930
rect -122 13903 216 13930
rect 268 13903 281 13955
rect 333 13903 347 13955
rect 399 13903 413 13955
rect 465 13903 479 13955
rect 531 13903 545 13955
rect 597 13903 611 13955
rect 663 13903 677 13955
rect 729 13903 887 13955
rect 939 13903 961 13955
rect 1013 13903 1035 13955
rect 1087 13903 1088 13955
rect -122 13881 1088 13903
rect -122 13878 216 13881
rect -778 13833 216 13878
rect -778 13829 -310 13833
rect -830 13807 -310 13829
rect -778 13781 -310 13807
rect -258 13781 -242 13833
rect -190 13781 -174 13833
rect -122 13829 216 13833
rect 268 13829 281 13881
rect 333 13829 347 13881
rect 399 13829 413 13881
rect 465 13829 479 13881
rect 531 13829 545 13881
rect 597 13829 611 13881
rect 663 13829 677 13881
rect 729 13829 887 13881
rect 939 13829 961 13881
rect 1013 13829 1035 13881
rect 1087 13829 1088 13881
rect -122 13807 1088 13829
rect -122 13781 216 13807
rect -778 13755 216 13781
rect 268 13755 281 13807
rect 333 13755 347 13807
rect 399 13755 413 13807
rect 465 13755 479 13807
rect 531 13755 545 13807
rect 597 13755 611 13807
rect 663 13755 677 13807
rect 729 13755 887 13807
rect 939 13755 961 13807
rect 1013 13755 1035 13807
rect 1087 13755 1088 13807
rect -830 13735 1088 13755
rect -830 13733 -310 13735
rect -778 13683 -310 13733
rect -258 13683 -242 13735
rect -190 13683 -174 13735
rect -122 13733 1088 13735
rect -122 13683 216 13733
rect -778 13681 216 13683
rect 268 13681 281 13733
rect 333 13681 347 13733
rect 399 13681 413 13733
rect 465 13681 479 13733
rect 531 13681 545 13733
rect 597 13681 611 13733
rect 663 13681 677 13733
rect 729 13681 887 13733
rect 939 13681 961 13733
rect 1013 13681 1035 13733
rect 1087 13681 1088 13733
rect -830 13675 1088 13681
rect -311 12114 -305 12166
rect -253 12114 -240 12166
rect -188 12114 -175 12166
rect -123 12114 -62 12166
rect -10 12114 8 12166
rect 60 12114 78 12166
rect 130 12114 148 12166
rect 200 12114 218 12166
rect 270 12114 289 12166
rect 341 12114 347 12166
rect -311 6391 -16 6397
rect -311 6339 -310 6391
rect -258 6339 -240 6391
rect -188 6339 -170 6391
rect -118 6339 -68 6391
rect -311 6321 -16 6339
rect -311 6269 -310 6321
rect -258 6269 -240 6321
rect -188 6269 -170 6321
rect -118 6269 -68 6321
rect -311 6251 -16 6269
rect -311 6199 -310 6251
rect -258 6199 -240 6251
rect -188 6199 -170 6251
rect -118 6199 -68 6251
rect -311 6181 -16 6199
rect -311 6129 -310 6181
rect -258 6129 -240 6181
rect -188 6129 -170 6181
rect -118 6129 -68 6181
rect -311 6111 -16 6129
rect -311 6059 -310 6111
rect -258 6059 -240 6111
rect -188 6059 -170 6111
rect -118 6059 -68 6111
rect -311 6041 -16 6059
rect -311 5989 -310 6041
rect -258 5989 -240 6041
rect -188 5989 -170 6041
rect -118 5989 -68 6041
rect -311 5971 -16 5989
rect -311 5919 -310 5971
rect -258 5919 -240 5971
rect -188 5919 -170 5971
rect -118 5919 -68 5971
rect -311 5901 -16 5919
rect -311 5849 -310 5901
rect -258 5849 -240 5901
rect -188 5849 -170 5901
rect -118 5849 -68 5901
rect -311 5830 -16 5849
rect -311 5778 -310 5830
rect -258 5778 -240 5830
rect -188 5778 -170 5830
rect -118 5778 -68 5830
rect -311 5772 -16 5778
rect -311 5070 -16 5076
rect -311 5018 -310 5070
rect -258 5018 -240 5070
rect -188 5018 -170 5070
rect -118 5018 -68 5070
rect -311 5004 -16 5018
rect -311 4952 -310 5004
rect -258 4952 -240 5004
rect -188 4952 -170 5004
rect -118 4952 -68 5004
rect -311 4938 -16 4952
rect -311 4886 -310 4938
rect -258 4886 -240 4938
rect -188 4886 -170 4938
rect -118 4886 -68 4938
rect -311 4872 -16 4886
rect -311 4820 -310 4872
rect -258 4820 -240 4872
rect -188 4820 -170 4872
rect -118 4820 -68 4872
rect -311 4806 -16 4820
rect -311 4754 -310 4806
rect -258 4754 -240 4806
rect -188 4754 -170 4806
rect -118 4754 -68 4806
rect -311 4740 -16 4754
rect -311 4688 -310 4740
rect -258 4688 -240 4740
rect -188 4688 -170 4740
rect -118 4688 -68 4740
rect -311 4674 -16 4688
rect -311 4622 -310 4674
rect -258 4622 -240 4674
rect -188 4622 -170 4674
rect -118 4622 -68 4674
rect -311 4607 -16 4622
rect -311 4555 -310 4607
rect -258 4555 -240 4607
rect -188 4555 -170 4607
rect -118 4555 -68 4607
rect -311 4540 -16 4555
rect -311 4488 -310 4540
rect -258 4488 -240 4540
rect -188 4488 -170 4540
rect -118 4488 -68 4540
rect -311 4473 -16 4488
rect -311 4421 -310 4473
rect -258 4421 -240 4473
rect -188 4421 -170 4473
rect -118 4421 -68 4473
rect -311 4406 -16 4421
rect -311 4354 -310 4406
rect -258 4354 -240 4406
rect -188 4354 -170 4406
rect -118 4354 -68 4406
rect -311 4339 -16 4354
rect -311 4287 -310 4339
rect -258 4287 -240 4339
rect -188 4287 -170 4339
rect -118 4287 -68 4339
rect -311 4272 -16 4287
rect -311 4220 -310 4272
rect -258 4220 -240 4272
rect -188 4220 -170 4272
rect -118 4220 -68 4272
rect -311 4205 -16 4220
rect -311 4153 -310 4205
rect -258 4153 -240 4205
rect -188 4153 -170 4205
rect -118 4153 -68 4205
rect 148 4691 585 4699
rect 148 4639 162 4691
rect 214 4639 585 4691
rect 148 4625 585 4639
rect 148 4573 162 4625
rect 214 4573 585 4625
rect 148 4558 585 4573
rect 148 4506 162 4558
rect 214 4506 585 4558
rect 148 4491 585 4506
rect 148 4439 162 4491
rect 214 4439 585 4491
rect 148 4424 585 4439
rect 148 4372 162 4424
rect 214 4372 585 4424
rect 148 4357 585 4372
rect 148 4305 162 4357
rect 214 4305 585 4357
rect 148 4290 585 4305
rect 148 4238 162 4290
rect 214 4238 585 4290
rect 148 4223 585 4238
rect 148 4171 162 4223
rect 214 4171 585 4223
rect 148 4162 585 4171
rect -311 4138 -16 4153
rect -311 4086 -310 4138
rect -258 4086 -240 4138
rect -188 4086 -170 4138
rect -118 4086 -68 4138
rect -311 4071 -16 4086
rect -311 4019 -310 4071
rect -258 4019 -240 4071
rect -188 4019 -170 4071
rect -118 4019 -68 4071
rect -311 4013 -16 4019
rect -830 2001 387 2007
rect -778 1999 387 2001
tri 387 1999 395 2007 sw
rect -778 1949 395 1999
rect -830 1919 395 1949
rect -778 1867 395 1919
rect -830 1861 395 1867
tri 327 1793 395 1861 ne
tri 395 1793 601 1999 sw
tri 395 1587 601 1793 ne
tri 601 1587 807 1793 sw
tri 601 1535 653 1587 ne
rect 653 1535 892 1587
rect 944 1535 961 1587
rect 1013 1535 1030 1587
rect 1082 1535 1088 1587
tri 653 1493 695 1535 ne
rect 695 1493 1088 1535
tri 695 1441 747 1493 ne
rect 747 1441 892 1493
rect 944 1441 961 1493
rect 1013 1441 1030 1493
rect 1082 1441 1088 1493
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_0
timestamp 1633016201
transform 1 0 456 0 1 1384
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_1
timestamp 1633016201
transform 1 0 456 0 1 2503
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_2
timestamp 1633016201
transform 1 0 456 0 1 3624
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_0
timestamp 1633016201
transform 1 0 415 0 -1 3593
box -28 0 148 471
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_1
timestamp 1633016201
transform 1 0 415 0 -1 4714
box -28 0 148 471
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_2
timestamp 1633016201
transform 1 0 415 0 -1 2472
box -28 0 148 471
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_3
timestamp 1633016201
transform 1 0 415 0 1 362
box -28 0 148 471
<< labels >>
flabel metal1 s 468 2328 508 2458 0 FreeSans 200 0 0 0 PD_H
port 1 nsew
flabel metal1 s 364 1833 410 1963 0 FreeSans 200 0 0 0 PAD
port 2 nsew
flabel metal1 s 364 2758 409 2888 0 FreeSans 200 0 0 0 PAD
port 2 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 3888486
string GDS_START 3582566
<< end >>


VVDD      vpwr0 GND  1.8
VNB       VNB  GND  0
VVGND     VGND GND  0

VC0 clk0 VGND pulse 0 1.8 6.18n 1n 1n 48n 100n
VC1 clk1 VGND pulse 0 1.8 7.52n 1n 1n 48n 100n
VC2 clk2 VGND pulse 0 1.8 5.03n 1n 1n 48n 100n
VC3 clk3 VGND pulse 0 1.8 7.79n 1n 1n 48n 100n
VC4 clk4 VGND pulse 0 1.8 3.22n 1n 1n 48n 100n
VC5 clk5 VGND pulse 0 1.8 7.55n 1n 1n 48n 100n
VC6 clk6 VGND pulse 0 1.8 5.45n 1n 1n 48n 100n
VC7 clk7 VGND pulse 0 1.8 7.91n 1n 1n 48n 100n
VC8 clk8 VGND pulse 0 1.8 6.88n 1n 1n 48n 100n
VC9 clk9 VGND pulse 0 1.8 5.91n 1n 1n 48n 100n
VC10 clk10 VGND pulse 0 1.8 1.21n 1n 1n 48n 100n
VC11 clk11 VGND pulse 0 1.8 3.19n 1n 1n 48n 100n
VC12 clk12 VGND pulse 0 1.8 2.14n 1n 1n 48n 100n
VC13 clk13 VGND pulse 0 1.8 2.1n 1n 1n 48n 100n
VC14 clk14 VGND pulse 0 1.8 2.08n 1n 1n 48n 100n
VC15 clk15 VGND pulse 0 1.8 6.97n 1n 1n 48n 100n
VC16 clk16 VGND pulse 0 1.8 1.86n 1n 1n 48n 100n
VC17 clk17 VGND pulse 0 1.8 5.89n 1n 1n 48n 100n
VC18 clk18 VGND pulse 0 1.8 2.73n 1n 1n 48n 100n
VC19 clk19 VGND pulse 0 1.8 3.4n 1n 1n 48n 100n
VC20 clk20 VGND pulse 0 1.8 7.9n 1n 1n 48n 100n
VC21 clk21 VGND pulse 0 1.8 3.68n 1n 1n 48n 100n
VC22 clk22 VGND pulse 0 1.8 6.48n 1n 1n 48n 100n
VC23 clk23 VGND pulse 0 1.8 2.29n 1n 1n 48n 100n
VC24 clk24 VGND pulse 0 1.8 5.07n 1n 1n 48n 100n
VC25 clk25 VGND pulse 0 1.8 3.56n 1n 1n 48n 100n
VC26 clk26 VGND pulse 0 1.8 4.75n 1n 1n 48n 100n
VC27 clk27 VGND pulse 0 1.8 6.03n 1n 1n 48n 100n
VC28 clk28 VGND pulse 0 1.8 6.65n 1n 1n 48n 100n
VC29 clk29 VGND pulse 0 1.8 1.98n 1n 1n 48n 100n
VC30 clk30 VGND pulse 0 1.8 6.97n 1n 1n 48n 100n
VC31 clk31 VGND pulse 0 1.8 4.2n 1n 1n 48n 100n

x00 clk0 VGND VNB vpwr0 vpwr0 co0 sky130_fd_sc_hd__clkbuf_1
x01 clk1 VGND VNB vpwr0 vpwr0 co1 sky130_fd_sc_hd__clkbuf_1
x02 clk2 VGND VNB vpwr0 vpwr0 co2 sky130_fd_sc_hd__clkbuf_1
x03 clk3 VGND VNB vpwr0 vpwr0 co3 sky130_fd_sc_hd__clkbuf_1
x04 clk4 VGND VNB vpwr0 vpwr0 co4 sky130_fd_sc_hd__clkbuf_1
x05 clk5 VGND VNB vpwr0 vpwr0 co5 sky130_fd_sc_hd__clkbuf_1
x06 clk6 VGND VNB vpwr0 vpwr0 co6 sky130_fd_sc_hd__clkbuf_1
x07 clk7 VGND VNB vpwr0 vpwr0 co7 sky130_fd_sc_hd__clkbuf_1
x08 clk8 VGND VNB vpwr0 vpwr0 co8 sky130_fd_sc_hd__clkbuf_1
x09 clk9 VGND VNB vpwr0 vpwr0 co9 sky130_fd_sc_hd__clkbuf_1
x010 clk10 VGND VNB vpwr0 vpwr0 co10 sky130_fd_sc_hd__clkbuf_1
x011 clk11 VGND VNB vpwr0 vpwr0 co11 sky130_fd_sc_hd__clkbuf_1
x012 clk12 VGND VNB vpwr0 vpwr0 co12 sky130_fd_sc_hd__clkbuf_1
x013 clk13 VGND VNB vpwr0 vpwr0 co13 sky130_fd_sc_hd__clkbuf_1
x014 clk14 VGND VNB vpwr0 vpwr0 co14 sky130_fd_sc_hd__clkbuf_1
x015 clk15 VGND VNB vpwr0 vpwr0 co15 sky130_fd_sc_hd__clkbuf_1
x016 clk16 VGND VNB vpwr0 vpwr0 co16 sky130_fd_sc_hd__clkbuf_1
x017 clk17 VGND VNB vpwr0 vpwr0 co17 sky130_fd_sc_hd__clkbuf_1
x018 clk18 VGND VNB vpwr0 vpwr0 co18 sky130_fd_sc_hd__clkbuf_1
x019 clk19 VGND VNB vpwr0 vpwr0 co19 sky130_fd_sc_hd__clkbuf_1
x020 clk20 VGND VNB vpwr0 vpwr0 co20 sky130_fd_sc_hd__clkbuf_1
x021 clk21 VGND VNB vpwr0 vpwr0 co21 sky130_fd_sc_hd__clkbuf_1
x022 clk22 VGND VNB vpwr0 vpwr0 co22 sky130_fd_sc_hd__clkbuf_1
x023 clk23 VGND VNB vpwr0 vpwr0 co23 sky130_fd_sc_hd__clkbuf_1
x024 clk24 VGND VNB vpwr0 vpwr0 co24 sky130_fd_sc_hd__clkbuf_1
x025 clk25 VGND VNB vpwr0 vpwr0 co25 sky130_fd_sc_hd__clkbuf_1
x026 clk26 VGND VNB vpwr0 vpwr0 co26 sky130_fd_sc_hd__clkbuf_1
x027 clk27 VGND VNB vpwr0 vpwr0 co27 sky130_fd_sc_hd__clkbuf_1
x028 clk28 VGND VNB vpwr0 vpwr0 co28 sky130_fd_sc_hd__clkbuf_1
x029 clk29 VGND VNB vpwr0 vpwr0 co29 sky130_fd_sc_hd__clkbuf_1
x030 clk30 VGND VNB vpwr0 vpwr0 co30 sky130_fd_sc_hd__clkbuf_1
x031 clk31 VGND VNB vpwr0 vpwr0 co31 sky130_fd_sc_hd__clkbuf_1

R0 co0 co1 50
R1 co1 co2 50
R2 co2 co3 50
R3 co3 co4 50
R4 co4 co5 50
R5 co5 co6 50
R6 co6 co7 50
R7 co7 co8 50
R8 co8 co9 50
R9 co9 co10 50
R10 co10 co11 50
R11 co11 co12 50
R12 co12 co13 50
R13 co13 co14 50
R14 co14 co15 50
R15 co15 co16 50
R16 co16 co17 50
R17 co17 co18 50
R18 co18 co19 50
R19 co19 co20 50
R20 co20 co21 50
R21 co21 co22 50
R22 co22 co23 50
R23 co23 co24 50
R24 co24 co25 50
R25 co25 co26 50
R26 co26 co27 50
R27 co27 co28 50
R28 co28 co29 50
R29 co29 co30 50
R30 co30 co31 50
R31 co31 co32 50

x10 co1 VGND VNB vpwr0 vpwr0 ff0 sky130_fd_sc_hd__clkbuf_16
x11 co2 VGND VNB vpwr0 vpwr0 ff1 sky130_fd_sc_hd__clkbuf_16
x12 co3 VGND VNB vpwr0 vpwr0 ff2 sky130_fd_sc_hd__clkbuf_16
x13 co4 VGND VNB vpwr0 vpwr0 ff3 sky130_fd_sc_hd__clkbuf_16
x14 co5 VGND VNB vpwr0 vpwr0 ff4 sky130_fd_sc_hd__clkbuf_16
x15 co6 VGND VNB vpwr0 vpwr0 ff5 sky130_fd_sc_hd__clkbuf_16
x16 co7 VGND VNB vpwr0 vpwr0 ff6 sky130_fd_sc_hd__clkbuf_16
x17 co8 VGND VNB vpwr0 vpwr0 ff7 sky130_fd_sc_hd__clkbuf_16
x18 co9 VGND VNB vpwr0 vpwr0 ff8 sky130_fd_sc_hd__clkbuf_16
x19 co10 VGND VNB vpwr0 vpwr0 ff9 sky130_fd_sc_hd__clkbuf_16
x110 co11 VGND VNB vpwr0 vpwr0 ff10 sky130_fd_sc_hd__clkbuf_16
x111 co12 VGND VNB vpwr0 vpwr0 ff11 sky130_fd_sc_hd__clkbuf_16
x112 co13 VGND VNB vpwr0 vpwr0 ff12 sky130_fd_sc_hd__clkbuf_16
x113 co14 VGND VNB vpwr0 vpwr0 ff13 sky130_fd_sc_hd__clkbuf_16
x114 co15 VGND VNB vpwr0 vpwr0 ff14 sky130_fd_sc_hd__clkbuf_16
x115 co16 VGND VNB vpwr0 vpwr0 ff15 sky130_fd_sc_hd__clkbuf_16
x116 co17 VGND VNB vpwr0 vpwr0 ff16 sky130_fd_sc_hd__clkbuf_16
x117 co18 VGND VNB vpwr0 vpwr0 ff17 sky130_fd_sc_hd__clkbuf_16
x118 co19 VGND VNB vpwr0 vpwr0 ff18 sky130_fd_sc_hd__clkbuf_16
x119 co20 VGND VNB vpwr0 vpwr0 ff19 sky130_fd_sc_hd__clkbuf_16
x120 co21 VGND VNB vpwr0 vpwr0 ff20 sky130_fd_sc_hd__clkbuf_16
x121 co22 VGND VNB vpwr0 vpwr0 ff21 sky130_fd_sc_hd__clkbuf_16
x122 co23 VGND VNB vpwr0 vpwr0 ff22 sky130_fd_sc_hd__clkbuf_16
x123 co24 VGND VNB vpwr0 vpwr0 ff23 sky130_fd_sc_hd__clkbuf_16
x124 co25 VGND VNB vpwr0 vpwr0 ff24 sky130_fd_sc_hd__clkbuf_16
x125 co26 VGND VNB vpwr0 vpwr0 ff25 sky130_fd_sc_hd__clkbuf_16
x126 co27 VGND VNB vpwr0 vpwr0 ff26 sky130_fd_sc_hd__clkbuf_16
x127 co28 VGND VNB vpwr0 vpwr0 ff27 sky130_fd_sc_hd__clkbuf_16
x128 co29 VGND VNB vpwr0 vpwr0 ff28 sky130_fd_sc_hd__clkbuf_16
x129 co30 VGND VNB vpwr0 vpwr0 ff29 sky130_fd_sc_hd__clkbuf_16
x130 co31 VGND VNB vpwr0 vpwr0 ff30 sky130_fd_sc_hd__clkbuf_16
x131 co32 VGND VNB vpwr0 vpwr0 ff31 sky130_fd_sc_hd__clkbuf_16

.lib /ciic/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /ciic/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.save clk0
.save clk1
.save clk2
.save clk3
.save clk4
.save clk5
.save clk6
.save clk7
.save clk8
.save clk9
.save clk10
.save clk11
.save clk12
.save clk13
.save clk14
.save clk15
.save clk16
.save clk17
.save clk18
.save clk19
.save clk20
.save clk21
.save clk22
.save clk23
.save clk24
.save clk25
.save clk26
.save clk27
.save clk28
.save clk29
.save clk30
.save clk31

.save co0
.save co1
.save co2
.save co3
.save co4
.save co5
.save co6
.save co7
.save co8
.save co9
.save co10
.save co11
.save co12
.save co13
.save co14
.save co15
.save co16
.save co17
.save co18
.save co19
.save co20
.save co21
.save co22
.save co23
.save co24
.save co25
.save co26
.save co27
.save co28
.save co29
.save co30
.save co31
.save co32

.save ff0
.save ff1
.save ff2
.save ff3
.save ff4
.save ff5
.save ff6
.save ff7
.save ff8
.save ff9
.save ff10
.save ff11
.save ff12
.save ff13
.save ff14
.save ff15
.save ff16
.save ff17
.save ff18
.save ff19
.save ff20
.save ff21
.save ff22
.save ff23
.save ff24
.save ff25
.save ff26
.save ff27
.save ff28
.save ff29
.save ff30
.save ff31

.save vpwr0
.save vpwr1
.save vpwr2
.save vpwr3
.save vpwr4
.save vpwr5
.save vpwr6
.save vpwr7
.save vpwr8
.save vpwr9
.save vpwr10
.save vpwr11
.save vpwr12
.save vpwr13
.save vpwr14
.save vpwr15
.save vpwr16
.save vpwr17
.save vpwr18
.save vpwr19
.save vpwr20
.save vpwr21
.save vpwr22
.save vpwr23
.save vpwr24
.save vpwr25
.save vpwr26
.save vpwr27
.save vpwr28
.save vpwr29
.save vpwr30
.save vpwr31


.save all
.options savecurrents
.tran 0.2n 300n

.end

magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1210 -1268 1844 2129
<< nwell >>
rect 50 482 584 814
<< pwell >>
rect 90 267 544 403
rect 136 -8 540 78
<< mvnmos >>
rect 169 293 289 377
rect 345 293 465 377
<< mvpmos >>
rect 169 548 289 748
rect 345 548 465 748
<< mvndiff >>
rect 116 339 169 377
rect 116 305 124 339
rect 158 305 169 339
rect 116 293 169 305
rect 289 339 345 377
rect 289 305 300 339
rect 334 305 345 339
rect 289 293 345 305
rect 465 339 518 377
rect 465 305 476 339
rect 510 305 518 339
rect 465 293 518 305
<< mvpdiff >>
rect 116 730 169 748
rect 116 696 124 730
rect 158 696 169 730
rect 116 662 169 696
rect 116 628 124 662
rect 158 628 169 662
rect 116 594 169 628
rect 116 560 124 594
rect 158 560 169 594
rect 116 548 169 560
rect 289 730 345 748
rect 289 696 300 730
rect 334 696 345 730
rect 289 662 345 696
rect 289 628 300 662
rect 334 628 345 662
rect 289 594 345 628
rect 289 560 300 594
rect 334 560 345 594
rect 289 548 345 560
rect 465 730 518 748
rect 465 696 476 730
rect 510 696 518 730
rect 465 662 518 696
rect 465 628 476 662
rect 510 628 518 662
rect 465 594 518 628
rect 465 560 476 594
rect 510 560 518 594
rect 465 548 518 560
<< mvndiffc >>
rect 124 305 158 339
rect 300 305 334 339
rect 476 305 510 339
<< mvpdiffc >>
rect 124 696 158 730
rect 124 628 158 662
rect 124 560 158 594
rect 300 696 334 730
rect 300 628 334 662
rect 300 560 334 594
rect 476 696 510 730
rect 476 628 510 662
rect 476 560 510 594
<< psubdiff >>
rect 162 18 186 52
rect 220 18 276 52
rect 310 18 366 52
rect 400 18 456 52
rect 490 18 514 52
<< psubdiffcont >>
rect 186 18 220 52
rect 276 18 310 52
rect 366 18 400 52
rect 456 18 490 52
<< poly >>
rect 169 748 289 780
rect 345 748 465 780
rect 169 493 289 548
rect 345 493 465 548
rect 169 477 465 493
rect 169 443 185 477
rect 219 443 261 477
rect 295 443 338 477
rect 372 443 415 477
rect 449 443 465 477
rect 169 427 465 443
rect 169 377 289 427
rect 345 377 465 427
rect 169 261 289 293
rect 345 261 465 293
<< polycont >>
rect 185 443 219 477
rect 261 443 295 477
rect 338 443 372 477
rect 415 443 449 477
<< locali >>
rect 124 734 158 746
rect 124 662 158 696
rect 124 594 158 628
rect 124 544 158 560
rect 300 730 334 746
rect 300 662 334 696
rect 300 594 334 628
rect 300 544 334 556
rect 476 734 510 746
rect 476 662 510 696
rect 476 594 510 628
rect 476 544 510 560
rect 169 443 185 477
rect 219 443 261 477
rect 295 443 338 477
rect 372 443 415 477
rect 449 443 465 477
rect 124 339 158 343
rect 300 339 334 361
rect 476 339 510 343
rect 162 52 514 58
rect 162 18 186 52
rect 228 18 276 52
rect 312 18 363 52
rect 400 18 448 52
rect 490 18 514 52
rect 162 12 514 18
<< viali >>
rect 124 730 158 734
rect 124 700 158 730
rect 124 628 158 662
rect 300 628 334 662
rect 300 560 334 590
rect 300 556 334 560
rect 476 730 510 734
rect 476 700 510 730
rect 476 628 510 662
rect 124 343 158 377
rect 124 271 158 305
rect 300 361 334 395
rect 300 305 334 323
rect 300 289 334 305
rect 476 343 510 377
rect 476 271 510 305
rect 194 18 220 52
rect 220 18 228 52
rect 278 18 310 52
rect 310 18 312 52
rect 363 18 366 52
rect 366 18 397 52
rect 448 18 456 52
rect 456 18 482 52
<< metal1 >>
rect 118 734 164 869
rect 118 700 124 734
rect 158 700 164 734
rect 118 662 164 700
rect 470 734 516 869
rect 470 700 476 734
rect 510 700 516 734
rect 118 628 124 662
rect 158 628 164 662
rect 118 616 164 628
rect 289 662 346 674
rect 289 628 300 662
rect 334 628 346 662
rect 289 590 346 628
rect 470 662 516 700
rect 470 628 476 662
rect 510 628 516 662
rect 470 616 516 628
rect 289 556 300 590
rect 334 556 346 590
rect 289 395 346 556
rect 118 377 164 389
rect 118 343 124 377
rect 158 343 164 377
rect 118 305 164 343
rect 118 271 124 305
rect 158 271 164 305
rect 289 361 300 395
rect 334 361 346 395
rect 289 323 346 361
rect 289 289 300 323
rect 334 289 346 323
rect 289 277 346 289
rect 470 377 516 389
rect 470 343 476 377
rect 510 343 516 377
rect 470 305 516 343
rect 118 58 164 271
rect 470 271 476 305
rect 510 271 516 305
rect 470 58 516 271
rect 118 52 516 58
rect 118 18 194 52
rect 228 18 278 52
rect 312 18 363 52
rect 397 18 448 52
rect 482 18 516 52
rect 118 12 516 18
use sky130_fd_pr__pfet_01v8__example_55959141808470  sky130_fd_pr__pfet_01v8__example_55959141808470_0
timestamp 1633016201
transform 1 0 169 0 1 548
box -28 0 324 97
use sky130_fd_pr__nfet_01v8__example_55959141808499  sky130_fd_pr__nfet_01v8__example_55959141808499_0
timestamp 1633016201
transform 1 0 169 0 1 293
box -28 0 324 29
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48518720
string GDS_START 48515308
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016076
<< checkpaint >>
rect -1260 -1260 2620 2478
<< pwell >>
rect 547 874 568 923
<< poly >>
rect 0 1202 1360 1218
rect 0 1168 80 1202
rect 114 1168 148 1202
rect 182 1168 216 1202
rect 250 1168 284 1202
rect 318 1168 352 1202
rect 386 1168 420 1202
rect 454 1168 488 1202
rect 522 1168 556 1202
rect 590 1168 624 1202
rect 658 1168 702 1202
rect 736 1168 770 1202
rect 804 1168 838 1202
rect 872 1168 906 1202
rect 940 1168 974 1202
rect 1008 1168 1042 1202
rect 1076 1168 1110 1202
rect 1144 1168 1178 1202
rect 1212 1168 1246 1202
rect 1280 1168 1360 1202
rect 0 1136 1360 1168
rect 0 1102 16 1136
rect 50 1102 1310 1136
rect 1344 1102 1360 1136
rect 0 1068 1360 1102
rect 0 1034 16 1068
rect 50 1034 1310 1068
rect 1344 1034 1360 1068
rect 0 1000 1360 1034
rect 0 966 16 1000
rect 50 966 1310 1000
rect 1344 966 1360 1000
rect 0 932 1360 966
rect 0 898 16 932
rect 50 898 1310 932
rect 1344 898 1360 932
rect 0 864 1360 898
rect 0 830 16 864
rect 50 830 1310 864
rect 1344 830 1360 864
rect 0 796 1360 830
rect 0 762 16 796
rect 50 762 1310 796
rect 1344 762 1360 796
rect 0 728 1360 762
rect 0 694 16 728
rect 50 694 1310 728
rect 1344 694 1360 728
rect 0 660 1360 694
rect 0 626 16 660
rect 50 626 1310 660
rect 1344 626 1360 660
rect 0 592 1360 626
rect 0 558 16 592
rect 50 558 1310 592
rect 1344 558 1360 592
rect 0 524 1360 558
rect 0 490 16 524
rect 50 490 1310 524
rect 1344 490 1360 524
rect 0 456 1360 490
rect 0 422 16 456
rect 50 422 1310 456
rect 1344 422 1360 456
rect 0 388 1360 422
rect 0 354 16 388
rect 50 354 1310 388
rect 1344 354 1360 388
rect 0 320 1360 354
rect 0 286 16 320
rect 50 286 1310 320
rect 1344 286 1360 320
rect 0 252 1360 286
rect 0 218 16 252
rect 50 218 1310 252
rect 1344 218 1360 252
rect 0 184 1360 218
rect 0 150 16 184
rect 50 150 1310 184
rect 1344 150 1360 184
rect 0 116 1360 150
rect 0 82 16 116
rect 50 82 1310 116
rect 1344 82 1360 116
rect 0 50 1360 82
rect 0 16 80 50
rect 114 16 148 50
rect 182 16 216 50
rect 250 16 284 50
rect 318 16 352 50
rect 386 16 420 50
rect 454 16 488 50
rect 522 16 556 50
rect 590 16 624 50
rect 658 16 702 50
rect 736 16 770 50
rect 804 16 838 50
rect 872 16 906 50
rect 940 16 974 50
rect 1008 16 1042 50
rect 1076 16 1110 50
rect 1144 16 1178 50
rect 1212 16 1246 50
rect 1280 16 1360 50
rect 0 0 1360 16
<< polycont >>
rect 80 1168 114 1202
rect 148 1168 182 1202
rect 216 1168 250 1202
rect 284 1168 318 1202
rect 352 1168 386 1202
rect 420 1168 454 1202
rect 488 1168 522 1202
rect 556 1168 590 1202
rect 624 1168 658 1202
rect 702 1168 736 1202
rect 770 1168 804 1202
rect 838 1168 872 1202
rect 906 1168 940 1202
rect 974 1168 1008 1202
rect 1042 1168 1076 1202
rect 1110 1168 1144 1202
rect 1178 1168 1212 1202
rect 1246 1168 1280 1202
rect 16 1102 50 1136
rect 1310 1102 1344 1136
rect 16 1034 50 1068
rect 1310 1034 1344 1068
rect 16 966 50 1000
rect 1310 966 1344 1000
rect 16 898 50 932
rect 1310 898 1344 932
rect 16 830 50 864
rect 1310 830 1344 864
rect 16 762 50 796
rect 1310 762 1344 796
rect 16 694 50 728
rect 1310 694 1344 728
rect 16 626 50 660
rect 1310 626 1344 660
rect 16 558 50 592
rect 1310 558 1344 592
rect 16 490 50 524
rect 1310 490 1344 524
rect 16 422 50 456
rect 1310 422 1344 456
rect 16 354 50 388
rect 1310 354 1344 388
rect 16 286 50 320
rect 1310 286 1344 320
rect 16 218 50 252
rect 1310 218 1344 252
rect 16 150 50 184
rect 1310 150 1344 184
rect 16 82 50 116
rect 1310 82 1344 116
rect 80 16 114 50
rect 148 16 182 50
rect 216 16 250 50
rect 284 16 318 50
rect 352 16 386 50
rect 420 16 454 50
rect 488 16 522 50
rect 556 16 590 50
rect 624 16 658 50
rect 702 16 736 50
rect 770 16 804 50
rect 838 16 872 50
rect 906 16 940 50
rect 974 16 1008 50
rect 1042 16 1076 50
rect 1110 16 1144 50
rect 1178 16 1212 50
rect 1246 16 1280 50
<< locali >>
rect 0 1202 1360 1218
rect 0 1168 80 1202
rect 116 1168 148 1202
rect 188 1168 216 1202
rect 260 1168 284 1202
rect 332 1168 352 1202
rect 404 1168 420 1202
rect 476 1168 488 1202
rect 548 1168 556 1202
rect 620 1168 624 1202
rect 658 1168 663 1202
rect 697 1168 702 1202
rect 736 1168 740 1202
rect 804 1168 812 1202
rect 872 1168 884 1202
rect 940 1168 956 1202
rect 1008 1168 1028 1202
rect 1076 1168 1100 1202
rect 1144 1168 1172 1202
rect 1212 1168 1244 1202
rect 1280 1168 1360 1202
rect 0 1152 1360 1168
rect 0 1136 66 1152
rect 0 1096 16 1136
rect 50 1096 66 1136
rect 1294 1136 1360 1152
rect 0 1068 66 1096
rect 100 1080 1260 1118
rect 1294 1096 1310 1136
rect 1344 1096 1360 1136
rect 0 1024 16 1068
rect 50 1046 66 1068
rect 648 1058 712 1080
rect 50 1024 611 1046
rect 0 1012 611 1024
rect 648 1024 663 1058
rect 697 1024 712 1058
rect 1294 1068 1360 1096
rect 1294 1046 1310 1068
rect 0 1000 66 1012
rect 0 952 16 1000
rect 50 952 66 1000
rect 648 986 712 1024
rect 746 1024 1310 1046
rect 1344 1024 1360 1068
rect 746 1012 1360 1024
rect 648 978 663 986
rect 0 932 66 952
rect 100 952 663 978
rect 697 978 712 986
rect 1294 1000 1360 1012
rect 697 952 1260 978
rect 100 940 1260 952
rect 1294 952 1310 1000
rect 1344 952 1360 1000
rect 0 880 16 932
rect 50 906 66 932
rect 648 914 712 940
rect 50 880 611 906
rect 0 872 611 880
rect 648 880 663 914
rect 697 880 712 914
rect 1294 932 1360 952
rect 1294 906 1310 932
rect 0 864 66 872
rect 0 808 16 864
rect 50 808 66 864
rect 648 842 712 880
rect 746 880 1310 906
rect 1344 880 1360 932
rect 746 872 1360 880
rect 648 838 663 842
rect 0 796 66 808
rect 100 808 663 838
rect 697 838 712 842
rect 1294 864 1360 872
rect 697 808 1260 838
rect 100 800 1260 808
rect 1294 808 1310 864
rect 1344 808 1360 864
rect 0 736 16 796
rect 50 766 66 796
rect 648 770 712 800
rect 50 736 611 766
rect 0 732 611 736
rect 648 736 663 770
rect 697 736 712 770
rect 1294 796 1360 808
rect 1294 766 1310 796
rect 0 728 66 732
rect 0 664 16 728
rect 50 664 66 728
rect 648 698 712 736
rect 746 736 1310 766
rect 1344 736 1360 796
rect 746 732 1360 736
rect 1294 728 1360 732
rect 0 660 66 664
rect 100 664 663 698
rect 697 664 1260 698
rect 100 660 1260 664
rect 1294 664 1310 728
rect 1344 664 1360 728
rect 1294 660 1360 664
rect 0 558 16 660
rect 50 626 66 660
rect 648 626 712 660
rect 1294 626 1310 660
rect 50 592 611 626
rect 648 592 663 626
rect 697 592 712 626
rect 746 592 1310 626
rect 50 558 66 592
rect 648 558 712 592
rect 1294 558 1310 592
rect 1344 558 1360 660
rect 0 554 66 558
rect 0 490 16 554
rect 50 490 66 554
rect 100 554 1260 558
rect 100 520 663 554
rect 697 520 1260 554
rect 1294 554 1360 558
rect 0 486 66 490
rect 0 482 611 486
rect 0 422 16 482
rect 50 452 611 482
rect 648 482 712 520
rect 1294 490 1310 554
rect 1344 490 1360 554
rect 1294 486 1360 490
rect 50 422 66 452
rect 0 410 66 422
rect 648 448 663 482
rect 697 448 712 482
rect 746 482 1360 486
rect 746 452 1310 482
rect 648 418 712 448
rect 1294 422 1310 452
rect 1344 422 1360 482
rect 0 354 16 410
rect 50 354 66 410
rect 100 410 1260 418
rect 100 380 663 410
rect 0 346 66 354
rect 648 376 663 380
rect 697 380 1260 410
rect 1294 410 1360 422
rect 697 376 712 380
rect 0 338 611 346
rect 0 286 16 338
rect 50 312 611 338
rect 648 338 712 376
rect 1294 354 1310 410
rect 1344 354 1360 410
rect 1294 346 1360 354
rect 50 286 66 312
rect 0 266 66 286
rect 648 304 663 338
rect 697 304 712 338
rect 746 338 1360 346
rect 746 312 1310 338
rect 648 278 712 304
rect 1294 286 1310 312
rect 1344 286 1360 338
rect 0 218 16 266
rect 50 218 66 266
rect 100 266 1260 278
rect 100 240 663 266
rect 0 206 66 218
rect 648 232 663 240
rect 697 240 1260 266
rect 1294 266 1360 286
rect 697 232 712 240
rect 0 194 611 206
rect 0 150 16 194
rect 50 172 611 194
rect 648 194 712 232
rect 1294 218 1310 266
rect 1344 218 1360 266
rect 1294 206 1360 218
rect 50 150 66 172
rect 0 122 66 150
rect 648 160 663 194
rect 697 160 712 194
rect 746 194 1360 206
rect 746 172 1310 194
rect 648 138 712 160
rect 1294 150 1310 172
rect 1344 150 1360 194
rect 0 82 16 122
rect 50 82 66 122
rect 100 100 1260 138
rect 1294 122 1360 150
rect 0 66 66 82
rect 1294 82 1310 122
rect 1344 82 1360 122
rect 1294 66 1360 82
rect 0 50 1360 66
rect 0 16 80 50
rect 116 16 148 50
rect 188 16 216 50
rect 260 16 284 50
rect 332 16 352 50
rect 404 16 420 50
rect 476 16 488 50
rect 548 16 556 50
rect 620 16 624 50
rect 658 16 663 50
rect 697 16 702 50
rect 736 16 740 50
rect 804 16 812 50
rect 872 16 884 50
rect 940 16 956 50
rect 1008 16 1028 50
rect 1076 16 1100 50
rect 1144 16 1172 50
rect 1212 16 1244 50
rect 1280 16 1360 50
rect 0 0 1360 16
<< viali >>
rect 82 1168 114 1202
rect 114 1168 116 1202
rect 154 1168 182 1202
rect 182 1168 188 1202
rect 226 1168 250 1202
rect 250 1168 260 1202
rect 298 1168 318 1202
rect 318 1168 332 1202
rect 370 1168 386 1202
rect 386 1168 404 1202
rect 442 1168 454 1202
rect 454 1168 476 1202
rect 514 1168 522 1202
rect 522 1168 548 1202
rect 586 1168 590 1202
rect 590 1168 620 1202
rect 663 1168 697 1202
rect 740 1168 770 1202
rect 770 1168 774 1202
rect 812 1168 838 1202
rect 838 1168 846 1202
rect 884 1168 906 1202
rect 906 1168 918 1202
rect 956 1168 974 1202
rect 974 1168 990 1202
rect 1028 1168 1042 1202
rect 1042 1168 1062 1202
rect 1100 1168 1110 1202
rect 1110 1168 1134 1202
rect 1172 1168 1178 1202
rect 1178 1168 1206 1202
rect 1244 1168 1246 1202
rect 1246 1168 1278 1202
rect 16 1102 50 1130
rect 16 1096 50 1102
rect 1310 1102 1344 1130
rect 1310 1096 1344 1102
rect 16 1034 50 1058
rect 16 1024 50 1034
rect 663 1024 697 1058
rect 16 966 50 986
rect 16 952 50 966
rect 1310 1034 1344 1058
rect 1310 1024 1344 1034
rect 663 952 697 986
rect 1310 966 1344 986
rect 1310 952 1344 966
rect 16 898 50 914
rect 16 880 50 898
rect 663 880 697 914
rect 16 830 50 842
rect 16 808 50 830
rect 1310 898 1344 914
rect 1310 880 1344 898
rect 663 808 697 842
rect 1310 830 1344 842
rect 1310 808 1344 830
rect 16 762 50 770
rect 16 736 50 762
rect 663 736 697 770
rect 16 694 50 698
rect 16 664 50 694
rect 1310 762 1344 770
rect 1310 736 1344 762
rect 663 664 697 698
rect 1310 694 1344 698
rect 1310 664 1344 694
rect 16 592 50 626
rect 663 592 697 626
rect 1310 592 1344 626
rect 16 524 50 554
rect 16 520 50 524
rect 663 520 697 554
rect 16 456 50 482
rect 16 448 50 456
rect 1310 524 1344 554
rect 1310 520 1344 524
rect 663 448 697 482
rect 1310 456 1344 482
rect 1310 448 1344 456
rect 16 388 50 410
rect 16 376 50 388
rect 663 376 697 410
rect 16 320 50 338
rect 16 304 50 320
rect 1310 388 1344 410
rect 1310 376 1344 388
rect 663 304 697 338
rect 1310 320 1344 338
rect 1310 304 1344 320
rect 16 252 50 266
rect 16 232 50 252
rect 663 232 697 266
rect 16 184 50 194
rect 16 160 50 184
rect 1310 252 1344 266
rect 1310 232 1344 252
rect 663 160 697 194
rect 1310 184 1344 194
rect 1310 160 1344 184
rect 16 116 50 122
rect 16 88 50 116
rect 1310 116 1344 122
rect 1310 88 1344 116
rect 82 16 114 50
rect 114 16 116 50
rect 154 16 182 50
rect 182 16 188 50
rect 226 16 250 50
rect 250 16 260 50
rect 298 16 318 50
rect 318 16 332 50
rect 370 16 386 50
rect 386 16 404 50
rect 442 16 454 50
rect 454 16 476 50
rect 514 16 522 50
rect 522 16 548 50
rect 586 16 590 50
rect 590 16 620 50
rect 663 16 697 50
rect 740 16 770 50
rect 770 16 774 50
rect 812 16 838 50
rect 838 16 846 50
rect 884 16 906 50
rect 906 16 918 50
rect 956 16 974 50
rect 974 16 990 50
rect 1028 16 1042 50
rect 1042 16 1062 50
rect 1100 16 1110 50
rect 1110 16 1134 50
rect 1172 16 1178 50
rect 1178 16 1206 50
rect 1244 16 1246 50
rect 1246 16 1278 50
<< metal1 >>
rect 0 1211 1360 1218
rect 0 1159 73 1211
rect 125 1159 137 1211
rect 189 1159 201 1211
rect 253 1202 265 1211
rect 317 1202 329 1211
rect 381 1202 393 1211
rect 445 1202 457 1211
rect 509 1202 521 1211
rect 573 1202 787 1211
rect 839 1202 851 1211
rect 903 1202 915 1211
rect 967 1202 979 1211
rect 1031 1202 1043 1211
rect 1095 1202 1107 1211
rect 260 1168 265 1202
rect 509 1168 514 1202
rect 573 1168 586 1202
rect 620 1168 663 1202
rect 697 1168 740 1202
rect 774 1168 787 1202
rect 846 1168 851 1202
rect 1095 1168 1100 1202
rect 253 1159 265 1168
rect 317 1159 329 1168
rect 381 1159 393 1168
rect 445 1159 457 1168
rect 509 1159 521 1168
rect 573 1159 787 1168
rect 839 1159 851 1168
rect 903 1159 915 1168
rect 967 1159 979 1168
rect 1031 1159 1043 1168
rect 1095 1159 1107 1168
rect 1159 1159 1171 1211
rect 1223 1159 1235 1211
rect 1287 1159 1360 1211
rect 0 1152 1360 1159
rect 0 1147 66 1152
rect 0 1095 7 1147
rect 59 1095 66 1147
rect 0 1083 66 1095
rect 0 1031 7 1083
rect 59 1031 66 1083
rect 0 1024 16 1031
rect 50 1024 66 1031
rect 0 1019 66 1024
rect 0 967 7 1019
rect 59 967 66 1019
rect 0 955 16 967
rect 50 955 66 967
rect 0 903 7 955
rect 59 903 66 955
rect 0 891 16 903
rect 50 891 66 903
rect 0 839 7 891
rect 59 839 66 891
rect 0 827 16 839
rect 50 827 66 839
rect 0 775 7 827
rect 59 775 66 827
rect 0 770 66 775
rect 0 763 16 770
rect 50 763 66 770
rect 0 711 7 763
rect 59 711 66 763
rect 0 698 66 711
rect 0 664 16 698
rect 50 664 66 698
rect 0 626 66 664
rect 0 592 16 626
rect 50 592 66 626
rect 0 554 66 592
rect 0 520 16 554
rect 50 520 66 554
rect 0 507 66 520
rect 0 455 7 507
rect 59 455 66 507
rect 0 448 16 455
rect 50 448 66 455
rect 0 443 66 448
rect 0 391 7 443
rect 59 391 66 443
rect 0 379 16 391
rect 50 379 66 391
rect 0 327 7 379
rect 59 327 66 379
rect 0 315 16 327
rect 50 315 66 327
rect 0 263 7 315
rect 59 263 66 315
rect 0 251 16 263
rect 50 251 66 263
rect 0 199 7 251
rect 59 199 66 251
rect 0 194 66 199
rect 0 187 16 194
rect 50 187 66 194
rect 0 135 7 187
rect 59 135 66 187
rect 0 123 66 135
rect 0 71 7 123
rect 59 71 66 123
rect 94 641 122 1124
rect 150 669 178 1152
rect 206 641 234 1124
rect 262 669 290 1152
rect 318 641 346 1124
rect 374 669 402 1152
rect 430 641 458 1124
rect 486 669 514 1152
rect 542 641 570 1124
rect 598 669 626 1152
rect 654 1115 706 1124
rect 654 1058 706 1063
rect 654 1051 663 1058
rect 697 1051 706 1058
rect 654 987 706 999
rect 654 923 706 935
rect 654 859 706 871
rect 654 795 706 807
rect 654 736 663 743
rect 697 736 706 743
rect 654 731 706 736
rect 654 664 663 679
rect 697 664 706 679
rect 734 669 762 1152
rect 654 641 706 664
rect 790 641 818 1124
rect 846 669 874 1152
rect 902 641 930 1124
rect 958 669 986 1152
rect 1014 641 1042 1124
rect 1070 669 1098 1152
rect 1126 641 1154 1124
rect 1182 669 1210 1152
rect 1294 1147 1360 1152
rect 1238 641 1266 1124
rect 94 635 1266 641
rect 94 583 105 635
rect 157 583 169 635
rect 221 583 233 635
rect 285 583 297 635
rect 349 583 361 635
rect 413 583 425 635
rect 477 583 489 635
rect 541 583 553 635
rect 605 583 617 635
rect 669 626 691 635
rect 669 583 691 592
rect 743 583 755 635
rect 807 583 819 635
rect 871 583 883 635
rect 935 583 947 635
rect 999 583 1011 635
rect 1063 583 1075 635
rect 1127 583 1139 635
rect 1191 583 1203 635
rect 1255 583 1266 635
rect 94 577 1266 583
rect 94 94 122 577
rect 0 66 66 71
rect 150 66 178 549
rect 206 94 234 577
rect 262 66 290 549
rect 318 94 346 577
rect 374 66 402 549
rect 430 94 458 577
rect 486 66 514 549
rect 542 94 570 577
rect 654 554 706 577
rect 598 66 626 549
rect 654 539 663 554
rect 697 539 706 554
rect 654 482 706 487
rect 654 475 663 482
rect 697 475 706 482
rect 654 411 706 423
rect 654 347 706 359
rect 654 283 706 295
rect 654 219 706 231
rect 654 160 663 167
rect 697 160 706 167
rect 654 155 706 160
rect 654 94 706 103
rect 734 66 762 549
rect 790 94 818 577
rect 846 66 874 549
rect 902 94 930 577
rect 958 66 986 549
rect 1014 94 1042 577
rect 1070 66 1098 549
rect 1126 94 1154 577
rect 1182 66 1210 549
rect 1238 94 1266 577
rect 1294 1095 1301 1147
rect 1353 1095 1360 1147
rect 1294 1083 1360 1095
rect 1294 1031 1301 1083
rect 1353 1031 1360 1083
rect 1294 1024 1310 1031
rect 1344 1024 1360 1031
rect 1294 1019 1360 1024
rect 1294 967 1301 1019
rect 1353 967 1360 1019
rect 1294 955 1310 967
rect 1344 955 1360 967
rect 1294 903 1301 955
rect 1353 903 1360 955
rect 1294 891 1310 903
rect 1344 891 1360 903
rect 1294 839 1301 891
rect 1353 839 1360 891
rect 1294 827 1310 839
rect 1344 827 1360 839
rect 1294 775 1301 827
rect 1353 775 1360 827
rect 1294 770 1360 775
rect 1294 763 1310 770
rect 1344 763 1360 770
rect 1294 711 1301 763
rect 1353 711 1360 763
rect 1294 698 1360 711
rect 1294 664 1310 698
rect 1344 664 1360 698
rect 1294 626 1360 664
rect 1294 592 1310 626
rect 1344 592 1360 626
rect 1294 554 1360 592
rect 1294 520 1310 554
rect 1344 520 1360 554
rect 1294 507 1360 520
rect 1294 455 1301 507
rect 1353 455 1360 507
rect 1294 448 1310 455
rect 1344 448 1360 455
rect 1294 443 1360 448
rect 1294 391 1301 443
rect 1353 391 1360 443
rect 1294 379 1310 391
rect 1344 379 1360 391
rect 1294 327 1301 379
rect 1353 327 1360 379
rect 1294 315 1310 327
rect 1344 315 1360 327
rect 1294 263 1301 315
rect 1353 263 1360 315
rect 1294 251 1310 263
rect 1344 251 1360 263
rect 1294 199 1301 251
rect 1353 199 1360 251
rect 1294 194 1360 199
rect 1294 187 1310 194
rect 1344 187 1360 194
rect 1294 135 1301 187
rect 1353 135 1360 187
rect 1294 123 1360 135
rect 1294 71 1301 123
rect 1353 71 1360 123
rect 1294 66 1360 71
rect 0 59 1360 66
rect 0 7 73 59
rect 125 7 137 59
rect 189 7 201 59
rect 253 50 265 59
rect 317 50 329 59
rect 381 50 393 59
rect 445 50 457 59
rect 509 50 521 59
rect 573 50 787 59
rect 839 50 851 59
rect 903 50 915 59
rect 967 50 979 59
rect 1031 50 1043 59
rect 1095 50 1107 59
rect 260 16 265 50
rect 509 16 514 50
rect 573 16 586 50
rect 620 16 663 50
rect 697 16 740 50
rect 774 16 787 50
rect 846 16 851 50
rect 1095 16 1100 50
rect 253 7 265 16
rect 317 7 329 16
rect 381 7 393 16
rect 445 7 457 16
rect 509 7 521 16
rect 573 7 787 16
rect 839 7 851 16
rect 903 7 915 16
rect 967 7 979 16
rect 1031 7 1043 16
rect 1095 7 1107 16
rect 1159 7 1171 59
rect 1223 7 1235 59
rect 1287 7 1360 59
rect 0 0 1360 7
<< via1 >>
rect 73 1202 125 1211
rect 73 1168 82 1202
rect 82 1168 116 1202
rect 116 1168 125 1202
rect 73 1159 125 1168
rect 137 1202 189 1211
rect 137 1168 154 1202
rect 154 1168 188 1202
rect 188 1168 189 1202
rect 137 1159 189 1168
rect 201 1202 253 1211
rect 265 1202 317 1211
rect 329 1202 381 1211
rect 393 1202 445 1211
rect 457 1202 509 1211
rect 521 1202 573 1211
rect 787 1202 839 1211
rect 851 1202 903 1211
rect 915 1202 967 1211
rect 979 1202 1031 1211
rect 1043 1202 1095 1211
rect 1107 1202 1159 1211
rect 201 1168 226 1202
rect 226 1168 253 1202
rect 265 1168 298 1202
rect 298 1168 317 1202
rect 329 1168 332 1202
rect 332 1168 370 1202
rect 370 1168 381 1202
rect 393 1168 404 1202
rect 404 1168 442 1202
rect 442 1168 445 1202
rect 457 1168 476 1202
rect 476 1168 509 1202
rect 521 1168 548 1202
rect 548 1168 573 1202
rect 787 1168 812 1202
rect 812 1168 839 1202
rect 851 1168 884 1202
rect 884 1168 903 1202
rect 915 1168 918 1202
rect 918 1168 956 1202
rect 956 1168 967 1202
rect 979 1168 990 1202
rect 990 1168 1028 1202
rect 1028 1168 1031 1202
rect 1043 1168 1062 1202
rect 1062 1168 1095 1202
rect 1107 1168 1134 1202
rect 1134 1168 1159 1202
rect 201 1159 253 1168
rect 265 1159 317 1168
rect 329 1159 381 1168
rect 393 1159 445 1168
rect 457 1159 509 1168
rect 521 1159 573 1168
rect 787 1159 839 1168
rect 851 1159 903 1168
rect 915 1159 967 1168
rect 979 1159 1031 1168
rect 1043 1159 1095 1168
rect 1107 1159 1159 1168
rect 1171 1202 1223 1211
rect 1171 1168 1172 1202
rect 1172 1168 1206 1202
rect 1206 1168 1223 1202
rect 1171 1159 1223 1168
rect 1235 1202 1287 1211
rect 1235 1168 1244 1202
rect 1244 1168 1278 1202
rect 1278 1168 1287 1202
rect 1235 1159 1287 1168
rect 7 1130 59 1147
rect 7 1096 16 1130
rect 16 1096 50 1130
rect 50 1096 59 1130
rect 7 1095 59 1096
rect 7 1058 59 1083
rect 7 1031 16 1058
rect 16 1031 50 1058
rect 50 1031 59 1058
rect 7 986 59 1019
rect 7 967 16 986
rect 16 967 50 986
rect 50 967 59 986
rect 7 952 16 955
rect 16 952 50 955
rect 50 952 59 955
rect 7 914 59 952
rect 7 903 16 914
rect 16 903 50 914
rect 50 903 59 914
rect 7 880 16 891
rect 16 880 50 891
rect 50 880 59 891
rect 7 842 59 880
rect 7 839 16 842
rect 16 839 50 842
rect 50 839 59 842
rect 7 808 16 827
rect 16 808 50 827
rect 50 808 59 827
rect 7 775 59 808
rect 7 736 16 763
rect 16 736 50 763
rect 50 736 59 763
rect 7 711 59 736
rect 7 482 59 507
rect 7 455 16 482
rect 16 455 50 482
rect 50 455 59 482
rect 7 410 59 443
rect 7 391 16 410
rect 16 391 50 410
rect 50 391 59 410
rect 7 376 16 379
rect 16 376 50 379
rect 50 376 59 379
rect 7 338 59 376
rect 7 327 16 338
rect 16 327 50 338
rect 50 327 59 338
rect 7 304 16 315
rect 16 304 50 315
rect 50 304 59 315
rect 7 266 59 304
rect 7 263 16 266
rect 16 263 50 266
rect 50 263 59 266
rect 7 232 16 251
rect 16 232 50 251
rect 50 232 59 251
rect 7 199 59 232
rect 7 160 16 187
rect 16 160 50 187
rect 50 160 59 187
rect 7 135 59 160
rect 7 122 59 123
rect 7 88 16 122
rect 16 88 50 122
rect 50 88 59 122
rect 7 71 59 88
rect 654 1063 706 1115
rect 654 1024 663 1051
rect 663 1024 697 1051
rect 697 1024 706 1051
rect 654 999 706 1024
rect 654 986 706 987
rect 654 952 663 986
rect 663 952 697 986
rect 697 952 706 986
rect 654 935 706 952
rect 654 914 706 923
rect 654 880 663 914
rect 663 880 697 914
rect 697 880 706 914
rect 654 871 706 880
rect 654 842 706 859
rect 654 808 663 842
rect 663 808 697 842
rect 697 808 706 842
rect 654 807 706 808
rect 654 770 706 795
rect 654 743 663 770
rect 663 743 697 770
rect 697 743 706 770
rect 654 698 706 731
rect 654 679 663 698
rect 663 679 697 698
rect 697 679 706 698
rect 105 583 157 635
rect 169 583 221 635
rect 233 583 285 635
rect 297 583 349 635
rect 361 583 413 635
rect 425 583 477 635
rect 489 583 541 635
rect 553 583 605 635
rect 617 626 669 635
rect 691 626 743 635
rect 617 592 663 626
rect 663 592 669 626
rect 691 592 697 626
rect 697 592 743 626
rect 617 583 669 592
rect 691 583 743 592
rect 755 583 807 635
rect 819 583 871 635
rect 883 583 935 635
rect 947 583 999 635
rect 1011 583 1063 635
rect 1075 583 1127 635
rect 1139 583 1191 635
rect 1203 583 1255 635
rect 654 520 663 539
rect 663 520 697 539
rect 697 520 706 539
rect 654 487 706 520
rect 654 448 663 475
rect 663 448 697 475
rect 697 448 706 475
rect 654 423 706 448
rect 654 410 706 411
rect 654 376 663 410
rect 663 376 697 410
rect 697 376 706 410
rect 654 359 706 376
rect 654 338 706 347
rect 654 304 663 338
rect 663 304 697 338
rect 697 304 706 338
rect 654 295 706 304
rect 654 266 706 283
rect 654 232 663 266
rect 663 232 697 266
rect 697 232 706 266
rect 654 231 706 232
rect 654 194 706 219
rect 654 167 663 194
rect 663 167 697 194
rect 697 167 706 194
rect 654 103 706 155
rect 1301 1130 1353 1147
rect 1301 1096 1310 1130
rect 1310 1096 1344 1130
rect 1344 1096 1353 1130
rect 1301 1095 1353 1096
rect 1301 1058 1353 1083
rect 1301 1031 1310 1058
rect 1310 1031 1344 1058
rect 1344 1031 1353 1058
rect 1301 986 1353 1019
rect 1301 967 1310 986
rect 1310 967 1344 986
rect 1344 967 1353 986
rect 1301 952 1310 955
rect 1310 952 1344 955
rect 1344 952 1353 955
rect 1301 914 1353 952
rect 1301 903 1310 914
rect 1310 903 1344 914
rect 1344 903 1353 914
rect 1301 880 1310 891
rect 1310 880 1344 891
rect 1344 880 1353 891
rect 1301 842 1353 880
rect 1301 839 1310 842
rect 1310 839 1344 842
rect 1344 839 1353 842
rect 1301 808 1310 827
rect 1310 808 1344 827
rect 1344 808 1353 827
rect 1301 775 1353 808
rect 1301 736 1310 763
rect 1310 736 1344 763
rect 1344 736 1353 763
rect 1301 711 1353 736
rect 1301 482 1353 507
rect 1301 455 1310 482
rect 1310 455 1344 482
rect 1344 455 1353 482
rect 1301 410 1353 443
rect 1301 391 1310 410
rect 1310 391 1344 410
rect 1344 391 1353 410
rect 1301 376 1310 379
rect 1310 376 1344 379
rect 1344 376 1353 379
rect 1301 338 1353 376
rect 1301 327 1310 338
rect 1310 327 1344 338
rect 1344 327 1353 338
rect 1301 304 1310 315
rect 1310 304 1344 315
rect 1344 304 1353 315
rect 1301 266 1353 304
rect 1301 263 1310 266
rect 1310 263 1344 266
rect 1344 263 1353 266
rect 1301 232 1310 251
rect 1310 232 1344 251
rect 1344 232 1353 251
rect 1301 199 1353 232
rect 1301 160 1310 187
rect 1310 160 1344 187
rect 1344 160 1353 187
rect 1301 135 1353 160
rect 1301 122 1353 123
rect 1301 88 1310 122
rect 1310 88 1344 122
rect 1344 88 1353 122
rect 1301 71 1353 88
rect 73 50 125 59
rect 73 16 82 50
rect 82 16 116 50
rect 116 16 125 50
rect 73 7 125 16
rect 137 50 189 59
rect 137 16 154 50
rect 154 16 188 50
rect 188 16 189 50
rect 137 7 189 16
rect 201 50 253 59
rect 265 50 317 59
rect 329 50 381 59
rect 393 50 445 59
rect 457 50 509 59
rect 521 50 573 59
rect 787 50 839 59
rect 851 50 903 59
rect 915 50 967 59
rect 979 50 1031 59
rect 1043 50 1095 59
rect 1107 50 1159 59
rect 201 16 226 50
rect 226 16 253 50
rect 265 16 298 50
rect 298 16 317 50
rect 329 16 332 50
rect 332 16 370 50
rect 370 16 381 50
rect 393 16 404 50
rect 404 16 442 50
rect 442 16 445 50
rect 457 16 476 50
rect 476 16 509 50
rect 521 16 548 50
rect 548 16 573 50
rect 787 16 812 50
rect 812 16 839 50
rect 851 16 884 50
rect 884 16 903 50
rect 915 16 918 50
rect 918 16 956 50
rect 956 16 967 50
rect 979 16 990 50
rect 990 16 1028 50
rect 1028 16 1031 50
rect 1043 16 1062 50
rect 1062 16 1095 50
rect 1107 16 1134 50
rect 1134 16 1159 50
rect 201 7 253 16
rect 265 7 317 16
rect 329 7 381 16
rect 393 7 445 16
rect 457 7 509 16
rect 521 7 573 16
rect 787 7 839 16
rect 851 7 903 16
rect 915 7 967 16
rect 979 7 1031 16
rect 1043 7 1095 16
rect 1107 7 1159 16
rect 1171 50 1223 59
rect 1171 16 1172 50
rect 1172 16 1206 50
rect 1206 16 1223 50
rect 1171 7 1223 16
rect 1235 50 1287 59
rect 1235 16 1244 50
rect 1244 16 1278 50
rect 1278 16 1287 50
rect 1235 7 1287 16
<< metal2 >>
rect 0 1213 619 1218
rect 0 1211 88 1213
rect 144 1211 168 1213
rect 224 1211 248 1213
rect 304 1211 328 1213
rect 384 1211 408 1213
rect 464 1211 488 1213
rect 544 1211 619 1213
rect 0 1159 73 1211
rect 317 1159 328 1211
rect 384 1159 393 1211
rect 573 1159 619 1211
rect 0 1157 88 1159
rect 144 1157 168 1159
rect 224 1157 248 1159
rect 304 1157 328 1159
rect 384 1157 408 1159
rect 464 1157 488 1159
rect 544 1157 619 1159
rect 0 1152 619 1157
rect 0 1147 66 1152
rect 0 1138 7 1147
rect 59 1138 66 1147
rect 0 1082 5 1138
rect 61 1082 66 1138
rect 647 1124 713 1218
rect 741 1213 1360 1218
rect 741 1211 818 1213
rect 874 1211 898 1213
rect 954 1211 978 1213
rect 1034 1211 1058 1213
rect 1114 1211 1138 1213
rect 1194 1211 1218 1213
rect 1274 1211 1360 1213
rect 741 1159 787 1211
rect 967 1159 978 1211
rect 1034 1159 1043 1211
rect 1287 1159 1360 1211
rect 741 1157 818 1159
rect 874 1157 898 1159
rect 954 1157 978 1159
rect 1034 1157 1058 1159
rect 1114 1157 1138 1159
rect 1194 1157 1218 1159
rect 1274 1157 1360 1159
rect 741 1152 1360 1157
rect 1294 1147 1360 1152
rect 1294 1138 1301 1147
rect 1353 1138 1360 1147
rect 94 1115 1266 1124
rect 94 1096 654 1115
rect 0 1058 7 1082
rect 59 1068 66 1082
rect 647 1077 654 1096
rect 706 1096 1266 1115
rect 706 1077 713 1096
rect 59 1058 619 1068
rect 0 1002 5 1058
rect 61 1040 619 1058
rect 61 1002 66 1040
rect 647 1021 651 1077
rect 707 1021 713 1077
rect 1294 1082 1299 1138
rect 1355 1082 1360 1138
rect 1294 1068 1301 1082
rect 741 1058 1301 1068
rect 1353 1058 1360 1082
rect 741 1040 1299 1058
rect 647 1012 654 1021
rect 0 978 7 1002
rect 59 978 66 1002
rect 94 999 654 1012
rect 706 1012 713 1021
rect 706 999 1266 1012
rect 94 997 1266 999
rect 94 984 651 997
rect 0 922 5 978
rect 61 956 66 978
rect 61 928 619 956
rect 647 941 651 984
rect 707 984 1266 997
rect 1294 1002 1299 1040
rect 1355 1002 1360 1058
rect 707 941 713 984
rect 1294 978 1301 1002
rect 1353 978 1360 1002
rect 1294 956 1299 978
rect 647 935 654 941
rect 706 935 713 941
rect 61 922 66 928
rect 0 903 7 922
rect 59 903 66 922
rect 0 898 66 903
rect 647 923 713 935
rect 741 928 1299 956
rect 647 917 654 923
rect 706 917 713 923
rect 647 900 651 917
rect 0 842 5 898
rect 61 844 66 898
rect 94 872 651 900
rect 647 861 651 872
rect 707 900 713 917
rect 1294 922 1299 928
rect 1355 922 1360 978
rect 1294 903 1301 922
rect 1353 903 1360 922
rect 707 872 1266 900
rect 1294 898 1360 903
rect 707 861 713 872
rect 647 859 713 861
rect 61 842 619 844
rect 0 839 7 842
rect 59 839 619 842
rect 0 827 619 839
rect 0 818 7 827
rect 59 818 619 827
rect 0 762 5 818
rect 61 816 619 818
rect 647 837 654 859
rect 706 837 713 859
rect 1294 844 1299 898
rect 61 762 66 816
rect 647 788 651 837
rect 0 738 7 762
rect 59 738 66 762
rect 94 781 651 788
rect 707 788 713 837
rect 741 842 1299 844
rect 1355 842 1360 898
rect 741 839 1301 842
rect 1353 839 1360 842
rect 741 827 1360 839
rect 741 818 1301 827
rect 1353 818 1360 827
rect 741 816 1299 818
rect 707 781 1266 788
rect 94 760 654 781
rect 0 682 5 738
rect 61 732 66 738
rect 647 757 654 760
rect 706 760 1266 781
rect 1294 762 1299 816
rect 1355 762 1360 818
rect 706 757 713 760
rect 61 682 619 732
rect 0 665 619 682
rect 647 701 651 757
rect 707 701 713 757
rect 1294 738 1301 762
rect 1353 738 1360 762
rect 1294 732 1299 738
rect 647 679 654 701
rect 706 679 713 701
rect 647 637 713 679
rect 741 682 1299 732
rect 1355 682 1360 738
rect 741 665 1360 682
rect 0 635 167 637
rect 223 635 247 637
rect 303 635 327 637
rect 383 635 407 637
rect 463 635 487 637
rect 543 635 567 637
rect 623 635 652 637
rect 708 635 737 637
rect 793 635 817 637
rect 873 635 897 637
rect 953 635 977 637
rect 1033 635 1057 637
rect 1113 635 1137 637
rect 1193 635 1360 637
rect 0 583 105 635
rect 157 583 167 635
rect 223 583 233 635
rect 477 583 487 635
rect 543 583 553 635
rect 807 583 817 635
rect 873 583 883 635
rect 1127 583 1137 635
rect 1193 583 1203 635
rect 1255 583 1360 635
rect 0 581 167 583
rect 223 581 247 583
rect 303 581 327 583
rect 383 581 407 583
rect 463 581 487 583
rect 543 581 567 583
rect 623 581 652 583
rect 708 581 737 583
rect 793 581 817 583
rect 873 581 897 583
rect 953 581 977 583
rect 1033 581 1057 583
rect 1113 581 1137 583
rect 1193 581 1360 583
rect 0 536 619 553
rect 0 480 5 536
rect 61 486 619 536
rect 647 539 713 581
rect 647 517 654 539
rect 706 517 713 539
rect 61 480 66 486
rect 0 456 7 480
rect 59 456 66 480
rect 647 461 651 517
rect 707 461 713 517
rect 741 536 1360 553
rect 741 486 1299 536
rect 647 458 654 461
rect 0 400 5 456
rect 61 402 66 456
rect 94 437 654 458
rect 706 458 713 461
rect 1294 480 1299 486
rect 1355 480 1360 536
rect 706 437 1266 458
rect 94 430 651 437
rect 61 400 619 402
rect 0 391 7 400
rect 59 391 619 400
rect 0 379 619 391
rect 0 376 7 379
rect 59 376 619 379
rect 0 320 5 376
rect 61 374 619 376
rect 647 381 651 430
rect 707 430 1266 437
rect 1294 456 1301 480
rect 1353 456 1360 480
rect 707 381 713 430
rect 1294 402 1299 456
rect 61 320 66 374
rect 647 359 654 381
rect 706 359 713 381
rect 741 400 1299 402
rect 1355 400 1360 456
rect 741 391 1301 400
rect 1353 391 1360 400
rect 741 379 1360 391
rect 741 376 1301 379
rect 1353 376 1360 379
rect 741 374 1299 376
rect 647 357 713 359
rect 647 346 651 357
rect 0 315 66 320
rect 94 318 651 346
rect 0 296 7 315
rect 59 296 66 315
rect 0 240 5 296
rect 61 290 66 296
rect 647 301 651 318
rect 707 346 713 357
rect 707 318 1266 346
rect 1294 320 1299 374
rect 1355 320 1360 376
rect 707 301 713 318
rect 647 295 654 301
rect 706 295 713 301
rect 61 262 619 290
rect 647 283 713 295
rect 1294 315 1360 320
rect 1294 296 1301 315
rect 1353 296 1360 315
rect 1294 290 1299 296
rect 647 277 654 283
rect 706 277 713 283
rect 61 240 66 262
rect 0 216 7 240
rect 59 216 66 240
rect 647 234 651 277
rect 0 160 5 216
rect 61 178 66 216
rect 94 221 651 234
rect 707 234 713 277
rect 741 262 1299 290
rect 1294 240 1299 262
rect 1355 240 1360 296
rect 707 221 1266 234
rect 94 219 1266 221
rect 94 206 654 219
rect 647 197 654 206
rect 706 206 1266 219
rect 1294 216 1301 240
rect 1353 216 1360 240
rect 706 197 713 206
rect 61 160 619 178
rect 0 136 7 160
rect 59 150 619 160
rect 59 136 66 150
rect 0 80 5 136
rect 61 80 66 136
rect 647 141 651 197
rect 707 141 713 197
rect 1294 178 1299 216
rect 741 160 1299 178
rect 1355 160 1360 216
rect 741 150 1301 160
rect 647 122 654 141
rect 94 103 654 122
rect 706 122 713 141
rect 1294 136 1301 150
rect 1353 136 1360 160
rect 706 103 1266 122
rect 94 94 1266 103
rect 0 71 7 80
rect 59 71 66 80
rect 0 66 66 71
rect 0 61 619 66
rect 0 59 88 61
rect 144 59 168 61
rect 224 59 248 61
rect 304 59 328 61
rect 384 59 408 61
rect 464 59 488 61
rect 544 59 619 61
rect 0 7 73 59
rect 317 7 328 59
rect 384 7 393 59
rect 573 7 619 59
rect 0 5 88 7
rect 144 5 168 7
rect 224 5 248 7
rect 304 5 328 7
rect 384 5 408 7
rect 464 5 488 7
rect 544 5 619 7
rect 0 0 619 5
rect 647 0 713 94
rect 1294 80 1299 136
rect 1355 80 1360 136
rect 1294 71 1301 80
rect 1353 71 1360 80
rect 1294 66 1360 71
rect 741 61 1360 66
rect 741 59 818 61
rect 874 59 898 61
rect 954 59 978 61
rect 1034 59 1058 61
rect 1114 59 1138 61
rect 1194 59 1218 61
rect 1274 59 1360 61
rect 741 7 787 59
rect 967 7 978 59
rect 1034 7 1043 59
rect 1287 7 1360 59
rect 741 5 818 7
rect 874 5 898 7
rect 954 5 978 7
rect 1034 5 1058 7
rect 1114 5 1138 7
rect 1194 5 1218 7
rect 1274 5 1360 7
rect 741 0 1360 5
<< via2 >>
rect 88 1211 144 1213
rect 168 1211 224 1213
rect 248 1211 304 1213
rect 328 1211 384 1213
rect 408 1211 464 1213
rect 488 1211 544 1213
rect 88 1159 125 1211
rect 125 1159 137 1211
rect 137 1159 144 1211
rect 168 1159 189 1211
rect 189 1159 201 1211
rect 201 1159 224 1211
rect 248 1159 253 1211
rect 253 1159 265 1211
rect 265 1159 304 1211
rect 328 1159 329 1211
rect 329 1159 381 1211
rect 381 1159 384 1211
rect 408 1159 445 1211
rect 445 1159 457 1211
rect 457 1159 464 1211
rect 488 1159 509 1211
rect 509 1159 521 1211
rect 521 1159 544 1211
rect 88 1157 144 1159
rect 168 1157 224 1159
rect 248 1157 304 1159
rect 328 1157 384 1159
rect 408 1157 464 1159
rect 488 1157 544 1159
rect 5 1095 7 1138
rect 7 1095 59 1138
rect 59 1095 61 1138
rect 5 1083 61 1095
rect 5 1082 7 1083
rect 7 1082 59 1083
rect 59 1082 61 1083
rect 818 1211 874 1213
rect 898 1211 954 1213
rect 978 1211 1034 1213
rect 1058 1211 1114 1213
rect 1138 1211 1194 1213
rect 1218 1211 1274 1213
rect 818 1159 839 1211
rect 839 1159 851 1211
rect 851 1159 874 1211
rect 898 1159 903 1211
rect 903 1159 915 1211
rect 915 1159 954 1211
rect 978 1159 979 1211
rect 979 1159 1031 1211
rect 1031 1159 1034 1211
rect 1058 1159 1095 1211
rect 1095 1159 1107 1211
rect 1107 1159 1114 1211
rect 1138 1159 1159 1211
rect 1159 1159 1171 1211
rect 1171 1159 1194 1211
rect 1218 1159 1223 1211
rect 1223 1159 1235 1211
rect 1235 1159 1274 1211
rect 818 1157 874 1159
rect 898 1157 954 1159
rect 978 1157 1034 1159
rect 1058 1157 1114 1159
rect 1138 1157 1194 1159
rect 1218 1157 1274 1159
rect 5 1031 7 1058
rect 7 1031 59 1058
rect 59 1031 61 1058
rect 5 1019 61 1031
rect 5 1002 7 1019
rect 7 1002 59 1019
rect 59 1002 61 1019
rect 651 1063 654 1077
rect 654 1063 706 1077
rect 706 1063 707 1077
rect 651 1051 707 1063
rect 651 1021 654 1051
rect 654 1021 706 1051
rect 706 1021 707 1051
rect 1299 1095 1301 1138
rect 1301 1095 1353 1138
rect 1353 1095 1355 1138
rect 1299 1083 1355 1095
rect 1299 1082 1301 1083
rect 1301 1082 1353 1083
rect 1353 1082 1355 1083
rect 651 987 707 997
rect 5 967 7 978
rect 7 967 59 978
rect 59 967 61 978
rect 5 955 61 967
rect 5 922 7 955
rect 7 922 59 955
rect 59 922 61 955
rect 651 941 654 987
rect 654 941 706 987
rect 706 941 707 987
rect 1299 1031 1301 1058
rect 1301 1031 1353 1058
rect 1353 1031 1355 1058
rect 1299 1019 1355 1031
rect 1299 1002 1301 1019
rect 1301 1002 1353 1019
rect 1353 1002 1355 1019
rect 1299 967 1301 978
rect 1301 967 1353 978
rect 1353 967 1355 978
rect 1299 955 1355 967
rect 5 891 61 898
rect 5 842 7 891
rect 7 842 59 891
rect 59 842 61 891
rect 651 871 654 917
rect 654 871 706 917
rect 706 871 707 917
rect 1299 922 1301 955
rect 1301 922 1353 955
rect 1353 922 1355 955
rect 651 861 707 871
rect 5 775 7 818
rect 7 775 59 818
rect 59 775 61 818
rect 1299 891 1355 898
rect 5 763 61 775
rect 5 762 7 763
rect 7 762 59 763
rect 59 762 61 763
rect 651 807 654 837
rect 654 807 706 837
rect 706 807 707 837
rect 651 795 707 807
rect 651 781 654 795
rect 654 781 706 795
rect 706 781 707 795
rect 1299 842 1301 891
rect 1301 842 1353 891
rect 1353 842 1355 891
rect 5 711 7 738
rect 7 711 59 738
rect 59 711 61 738
rect 1299 775 1301 818
rect 1301 775 1353 818
rect 1353 775 1355 818
rect 1299 763 1355 775
rect 1299 762 1301 763
rect 1301 762 1353 763
rect 1353 762 1355 763
rect 5 682 61 711
rect 651 743 654 757
rect 654 743 706 757
rect 706 743 707 757
rect 651 731 707 743
rect 651 701 654 731
rect 654 701 706 731
rect 706 701 707 731
rect 1299 711 1301 738
rect 1301 711 1353 738
rect 1353 711 1355 738
rect 1299 682 1355 711
rect 167 635 223 637
rect 247 635 303 637
rect 327 635 383 637
rect 407 635 463 637
rect 487 635 543 637
rect 567 635 623 637
rect 652 635 708 637
rect 737 635 793 637
rect 817 635 873 637
rect 897 635 953 637
rect 977 635 1033 637
rect 1057 635 1113 637
rect 1137 635 1193 637
rect 167 583 169 635
rect 169 583 221 635
rect 221 583 223 635
rect 247 583 285 635
rect 285 583 297 635
rect 297 583 303 635
rect 327 583 349 635
rect 349 583 361 635
rect 361 583 383 635
rect 407 583 413 635
rect 413 583 425 635
rect 425 583 463 635
rect 487 583 489 635
rect 489 583 541 635
rect 541 583 543 635
rect 567 583 605 635
rect 605 583 617 635
rect 617 583 623 635
rect 652 583 669 635
rect 669 583 691 635
rect 691 583 708 635
rect 737 583 743 635
rect 743 583 755 635
rect 755 583 793 635
rect 817 583 819 635
rect 819 583 871 635
rect 871 583 873 635
rect 897 583 935 635
rect 935 583 947 635
rect 947 583 953 635
rect 977 583 999 635
rect 999 583 1011 635
rect 1011 583 1033 635
rect 1057 583 1063 635
rect 1063 583 1075 635
rect 1075 583 1113 635
rect 1137 583 1139 635
rect 1139 583 1191 635
rect 1191 583 1193 635
rect 167 581 223 583
rect 247 581 303 583
rect 327 581 383 583
rect 407 581 463 583
rect 487 581 543 583
rect 567 581 623 583
rect 652 581 708 583
rect 737 581 793 583
rect 817 581 873 583
rect 897 581 953 583
rect 977 581 1033 583
rect 1057 581 1113 583
rect 1137 581 1193 583
rect 5 507 61 536
rect 5 480 7 507
rect 7 480 59 507
rect 59 480 61 507
rect 651 487 654 517
rect 654 487 706 517
rect 706 487 707 517
rect 651 475 707 487
rect 651 461 654 475
rect 654 461 706 475
rect 706 461 707 475
rect 1299 507 1355 536
rect 5 455 7 456
rect 7 455 59 456
rect 59 455 61 456
rect 5 443 61 455
rect 5 400 7 443
rect 7 400 59 443
rect 59 400 61 443
rect 1299 480 1301 507
rect 1301 480 1353 507
rect 1353 480 1355 507
rect 5 327 7 376
rect 7 327 59 376
rect 59 327 61 376
rect 651 423 654 437
rect 654 423 706 437
rect 706 423 707 437
rect 651 411 707 423
rect 651 381 654 411
rect 654 381 706 411
rect 706 381 707 411
rect 1299 455 1301 456
rect 1301 455 1353 456
rect 1353 455 1355 456
rect 1299 443 1355 455
rect 5 320 61 327
rect 1299 400 1301 443
rect 1301 400 1353 443
rect 1353 400 1355 443
rect 651 347 707 357
rect 5 263 7 296
rect 7 263 59 296
rect 59 263 61 296
rect 651 301 654 347
rect 654 301 706 347
rect 706 301 707 347
rect 1299 327 1301 376
rect 1301 327 1353 376
rect 1353 327 1355 376
rect 1299 320 1355 327
rect 5 251 61 263
rect 5 240 7 251
rect 7 240 59 251
rect 59 240 61 251
rect 5 199 7 216
rect 7 199 59 216
rect 59 199 61 216
rect 5 187 61 199
rect 5 160 7 187
rect 7 160 59 187
rect 59 160 61 187
rect 651 231 654 277
rect 654 231 706 277
rect 706 231 707 277
rect 1299 263 1301 296
rect 1301 263 1353 296
rect 1353 263 1355 296
rect 1299 251 1355 263
rect 1299 240 1301 251
rect 1301 240 1353 251
rect 1353 240 1355 251
rect 651 221 707 231
rect 5 135 7 136
rect 7 135 59 136
rect 59 135 61 136
rect 5 123 61 135
rect 5 80 7 123
rect 7 80 59 123
rect 59 80 61 123
rect 651 167 654 197
rect 654 167 706 197
rect 706 167 707 197
rect 651 155 707 167
rect 651 141 654 155
rect 654 141 706 155
rect 706 141 707 155
rect 1299 199 1301 216
rect 1301 199 1353 216
rect 1353 199 1355 216
rect 1299 187 1355 199
rect 1299 160 1301 187
rect 1301 160 1353 187
rect 1353 160 1355 187
rect 88 59 144 61
rect 168 59 224 61
rect 248 59 304 61
rect 328 59 384 61
rect 408 59 464 61
rect 488 59 544 61
rect 88 7 125 59
rect 125 7 137 59
rect 137 7 144 59
rect 168 7 189 59
rect 189 7 201 59
rect 201 7 224 59
rect 248 7 253 59
rect 253 7 265 59
rect 265 7 304 59
rect 328 7 329 59
rect 329 7 381 59
rect 381 7 384 59
rect 408 7 445 59
rect 445 7 457 59
rect 457 7 464 59
rect 488 7 509 59
rect 509 7 521 59
rect 521 7 544 59
rect 88 5 144 7
rect 168 5 224 7
rect 248 5 304 7
rect 328 5 384 7
rect 408 5 464 7
rect 488 5 544 7
rect 1299 135 1301 136
rect 1301 135 1353 136
rect 1353 135 1355 136
rect 1299 123 1355 135
rect 1299 80 1301 123
rect 1301 80 1353 123
rect 1353 80 1355 123
rect 818 59 874 61
rect 898 59 954 61
rect 978 59 1034 61
rect 1058 59 1114 61
rect 1138 59 1194 61
rect 1218 59 1274 61
rect 818 7 839 59
rect 839 7 851 59
rect 851 7 874 59
rect 898 7 903 59
rect 903 7 915 59
rect 915 7 954 59
rect 978 7 979 59
rect 979 7 1031 59
rect 1031 7 1034 59
rect 1058 7 1095 59
rect 1095 7 1107 59
rect 1107 7 1114 59
rect 1138 7 1159 59
rect 1159 7 1171 59
rect 1171 7 1194 59
rect 1218 7 1223 59
rect 1223 7 1235 59
rect 1235 7 1274 59
rect 818 5 874 7
rect 898 5 954 7
rect 978 5 1034 7
rect 1058 5 1114 7
rect 1138 5 1194 7
rect 1218 5 1274 7
<< metal3 >>
rect 0 1213 1360 1218
rect 0 1157 88 1213
rect 144 1157 168 1213
rect 224 1157 248 1213
rect 304 1157 328 1213
rect 384 1157 408 1213
rect 464 1157 488 1213
rect 544 1157 818 1213
rect 874 1157 898 1213
rect 954 1157 978 1213
rect 1034 1157 1058 1213
rect 1114 1157 1138 1213
rect 1194 1157 1218 1213
rect 1274 1157 1360 1213
rect 0 1152 1360 1157
rect 0 1138 66 1152
rect 0 1082 5 1138
rect 61 1082 66 1138
rect 0 1058 66 1082
rect 0 1002 5 1058
rect 61 1002 66 1058
rect 0 978 66 1002
rect 0 922 5 978
rect 61 922 66 978
rect 0 898 66 922
rect 0 842 5 898
rect 61 842 66 898
rect 0 818 66 842
rect 0 762 5 818
rect 61 762 66 818
rect 0 738 66 762
rect 0 682 5 738
rect 61 682 66 738
rect 0 536 66 682
rect 0 480 5 536
rect 61 480 66 536
rect 0 456 66 480
rect 0 400 5 456
rect 61 400 66 456
rect 0 376 66 400
rect 0 320 5 376
rect 61 320 66 376
rect 0 296 66 320
rect 0 240 5 296
rect 61 240 66 296
rect 0 216 66 240
rect 0 160 5 216
rect 61 160 66 216
rect 0 136 66 160
rect 0 80 5 136
rect 61 80 66 136
rect 126 642 194 1092
rect 254 702 322 1152
rect 382 642 450 1092
rect 510 702 578 1152
rect 638 1077 722 1092
rect 638 1021 651 1077
rect 707 1021 722 1077
rect 638 997 722 1021
rect 638 941 651 997
rect 707 941 722 997
rect 638 917 722 941
rect 638 861 651 917
rect 707 861 722 917
rect 638 837 722 861
rect 638 781 651 837
rect 707 781 722 837
rect 638 757 722 781
rect 638 701 651 757
rect 707 701 722 757
rect 782 702 850 1152
rect 638 642 722 701
rect 910 642 978 1092
rect 1038 702 1106 1152
rect 1294 1138 1360 1152
rect 1166 642 1234 1092
rect 126 637 1234 642
rect 126 581 167 637
rect 223 581 247 637
rect 303 581 327 637
rect 383 581 407 637
rect 463 581 487 637
rect 543 581 567 637
rect 623 581 652 637
rect 708 581 737 637
rect 793 581 817 637
rect 873 581 897 637
rect 953 581 977 637
rect 1033 581 1057 637
rect 1113 581 1137 637
rect 1193 581 1234 637
rect 126 576 1234 581
rect 126 126 194 576
rect 0 66 66 80
rect 254 66 322 516
rect 382 126 450 576
rect 638 517 722 576
rect 510 66 578 516
rect 638 461 651 517
rect 707 461 722 517
rect 638 437 722 461
rect 638 381 651 437
rect 707 381 722 437
rect 638 357 722 381
rect 638 301 651 357
rect 707 301 722 357
rect 638 277 722 301
rect 638 221 651 277
rect 707 221 722 277
rect 638 197 722 221
rect 638 141 651 197
rect 707 141 722 197
rect 638 126 722 141
rect 782 66 850 516
rect 910 126 978 576
rect 1038 66 1106 516
rect 1166 126 1234 576
rect 1294 1082 1299 1138
rect 1355 1082 1360 1138
rect 1294 1058 1360 1082
rect 1294 1002 1299 1058
rect 1355 1002 1360 1058
rect 1294 978 1360 1002
rect 1294 922 1299 978
rect 1355 922 1360 978
rect 1294 898 1360 922
rect 1294 842 1299 898
rect 1355 842 1360 898
rect 1294 818 1360 842
rect 1294 762 1299 818
rect 1355 762 1360 818
rect 1294 738 1360 762
rect 1294 682 1299 738
rect 1355 682 1360 738
rect 1294 536 1360 682
rect 1294 480 1299 536
rect 1355 480 1360 536
rect 1294 456 1360 480
rect 1294 400 1299 456
rect 1355 400 1360 456
rect 1294 376 1360 400
rect 1294 320 1299 376
rect 1355 320 1360 376
rect 1294 296 1360 320
rect 1294 240 1299 296
rect 1355 240 1360 296
rect 1294 216 1360 240
rect 1294 160 1299 216
rect 1355 160 1360 216
rect 1294 136 1360 160
rect 1294 80 1299 136
rect 1355 80 1360 136
rect 1294 66 1360 80
rect 0 61 1360 66
rect 0 5 88 61
rect 144 5 168 61
rect 224 5 248 61
rect 304 5 328 61
rect 384 5 408 61
rect 464 5 488 61
rect 544 5 818 61
rect 874 5 898 61
rect 954 5 978 61
rect 1034 5 1058 61
rect 1114 5 1138 61
rect 1194 5 1218 61
rect 1274 5 1360 61
rect 0 0 1360 5
<< metal4 >>
rect 0 0 1360 1218
<< comment >>
rect 617 1184 618 1218
rect 647 1216 713 1217
rect 34 34 1326 1184
<< labels >>
flabel metal4 s 788 902 841 957 3 FreeSans 520 0 0 0 MET4
port 3 nsew
flabel metal2 s 547 1174 566 1194 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 652 1169 704 1205 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 547 874 568 923 0 FreeSans 2000 0 0 0 SUB
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 187146
string GDS_START 160268
<< end >>

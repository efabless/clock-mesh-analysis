magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1288 -1260 1656 1357
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_0
timestamp 1633016201
transform 1 0 50 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_1
timestamp 1633016201
transform 1 0 156 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_2
timestamp 1633016201
transform 1 0 262 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1633016201
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_1
timestamp 1633016201
transform 1 0 368 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 396 97 396 97 0 FreeSans 300 0 0 0 S
flabel comment s 290 97 290 97 0 FreeSans 300 0 0 0 D
flabel comment s 184 97 184 97 0 FreeSans 300 0 0 0 S
flabel comment s 78 97 78 97 0 FreeSans 300 0 0 0 D
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 2233394
string GDS_START 2230978
<< end >>

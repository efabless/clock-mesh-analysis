magic
tech sky130A
magscale 1 2
timestamp 1633016214
<< metal4 >>
rect 0 13600 1000 18593
rect 0 12410 1000 13300
rect 0 11240 1000 12130
rect 0 10218 1000 10814
rect 0 9266 1000 9862
rect 0 7910 1000 8840
rect 0 5970 1000 6660
rect 0 4760 1000 5690
rect 0 3550 1000 4480
rect 0 1370 1000 2300
rect 0 0 1000 1090
<< obsm4 >>
rect 0 34750 1000 39593
<< metal5 >>
rect 0 34750 1000 39593
rect 0 13600 1000 18590
rect 0 12430 1000 13280
rect 0 11260 1000 12110
rect 0 7930 1000 8820
rect 0 5990 1000 6640
rect 0 4780 1000 5670
rect 0 3570 1000 4460
rect 0 1390 1000 2280
rect 0 20 1000 1070
<< labels >>
rlabel metal4 s 0 10218 1000 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 1000 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 0 5990 1000 6640 6 VSWITCH
port 3 nsew power bidirectional
rlabel metal4 s 0 5970 1000 6660 6 VSWITCH
port 3 nsew power bidirectional
rlabel metal5 s 0 12430 1000 13280 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal4 s 0 12410 1000 13300 6 VDDIO_Q
port 4 nsew power bidirectional
rlabel metal5 s 0 20 1000 1070 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal4 s 0 0 1000 1090 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal4 s 0 3550 1000 4480 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 0 13600 1000 18590 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 0 13600 1000 18593 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 0 3570 1000 4460 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 0 1390 1000 2280 6 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 0 1370 1000 2300 6 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 0 4780 1000 5670 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal4 s 0 4760 1000 5690 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal5 s 0 34750 1000 39593 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal5 s 0 7930 1000 8820 6 VSSD
port 9 nsew ground bidirectional
rlabel metal4 s 0 7910 1000 8840 6 VSSD
port 9 nsew ground bidirectional
rlabel metal5 s 0 11260 1000 12110 6 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal4 s 0 11240 1000 12130 6 VSSIO_Q
port 10 nsew ground bidirectional
<< properties >>
string LEFclass PAD AREAIO
string FIXED_BBOX 0 0 1000 39593
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__disconnect_vdda_slice_5um.gds
string GDS_END 7104
string GDS_START 170
<< end >>

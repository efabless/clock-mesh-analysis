magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1285 -1260 13309 1760
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_0
timestamp 1633016201
transform 1 0 641 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_1
timestamp 1633016201
transform 1 0 1633 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_2
timestamp 1633016201
transform 1 0 2625 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_3
timestamp 1633016201
transform 1 0 3617 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_4
timestamp 1633016201
transform 1 0 4609 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_5
timestamp 1633016201
transform 1 0 5601 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_6
timestamp 1633016201
transform 1 0 6593 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_7
timestamp 1633016201
transform 1 0 7585 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_8
timestamp 1633016201
transform 1 0 8577 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_9
timestamp 1633016201
transform 1 0 9569 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_10
timestamp 1633016201
transform 1 0 10561 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_11
timestamp 1633016201
transform 1 0 11553 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 12049 500 12049 500 0 FreeSans 300 0 0 0 D
flabel comment s 11683 481 11683 481 0 FreeSans 300 0 0 0 S
flabel comment s 11187 500 11187 500 0 FreeSans 300 0 0 0 D
flabel comment s 10691 481 10691 481 0 FreeSans 300 0 0 0 S
flabel comment s 10195 500 10195 500 0 FreeSans 300 0 0 0 D
flabel comment s 9699 481 9699 481 0 FreeSans 300 0 0 0 S
flabel comment s 9203 500 9203 500 0 FreeSans 300 0 0 0 D
flabel comment s 8707 481 8707 481 0 FreeSans 300 0 0 0 S
flabel comment s 8211 500 8211 500 0 FreeSans 300 0 0 0 D
flabel comment s 7715 481 7715 481 0 FreeSans 300 0 0 0 S
flabel comment s 7219 500 7219 500 0 FreeSans 300 0 0 0 D
flabel comment s 6723 481 6723 481 0 FreeSans 300 0 0 0 S
flabel comment s 6227 500 6227 500 0 FreeSans 300 0 0 0 D
flabel comment s 5731 481 5731 481 0 FreeSans 300 0 0 0 S
flabel comment s 5235 500 5235 500 0 FreeSans 300 0 0 0 D
flabel comment s 4739 481 4739 481 0 FreeSans 300 0 0 0 S
flabel comment s 4243 500 4243 500 0 FreeSans 300 0 0 0 D
flabel comment s 3747 481 3747 481 0 FreeSans 300 0 0 0 S
flabel comment s 3251 500 3251 500 0 FreeSans 300 0 0 0 D
flabel comment s 2755 481 2755 481 0 FreeSans 300 0 0 0 S
flabel comment s 2259 500 2259 500 0 FreeSans 300 0 0 0 D
flabel comment s 1763 481 1763 481 0 FreeSans 300 0 0 0 S
flabel comment s 1267 500 1267 500 0 FreeSans 300 0 0 0 D
flabel comment s 771 481 771 481 0 FreeSans 300 0 0 0 S
flabel comment s 275 500 275 500 0 FreeSans 300 0 0 0 D
flabel comment s -25 500 -25 500 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 3963174
string GDS_START 3950198
<< end >>


VVDD      vpwr_0 0  ${VDDD}
VNB       VNB  0  0
VVGND     VGND 0  0

RP_clk_buf1_0 vpwr_0 vpwr_clk_buf1_branch_0  ${R_clk_buf1_BASE}
RP_clk_buf1_1 vpwr_0 vpwr_clk_buf1_branch_1  ${R_clk_buf1_BASE}
RP_clk_buf1_2 vpwr_0 vpwr_clk_buf1_branch_2  ${R_clk_buf1_BASE}
RP_clk_buf1_3 vpwr_0 vpwr_clk_buf1_branch_3  ${R_clk_buf1_BASE}
RP_clk_buf1_4 vpwr_0 vpwr_clk_buf1_branch_4  ${R_clk_buf1_BASE}
RP_clk_buf1_5 vpwr_0 vpwr_clk_buf1_branch_5  ${R_clk_buf1_BASE}
RP_clk_buf1_6 vpwr_0 vpwr_clk_buf1_branch_6  ${R_clk_buf1_BASE}
RP_clk_buf1_LOAD_0  vpwr_clk_buf1_branch_0 vpwr_clk_buf1_0 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_1  vpwr_clk_buf1_branch_1 vpwr_clk_buf1_1 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_2  vpwr_clk_buf1_branch_2 vpwr_clk_buf1_2 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_3  vpwr_clk_buf1_branch_3 vpwr_clk_buf1_3 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_4  vpwr_clk_buf1_branch_4 vpwr_clk_buf1_4 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_5  vpwr_clk_buf1_branch_5 vpwr_clk_buf1_5 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_6  vpwr_clk_buf1_branch_6 vpwr_clk_buf1_6 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_7  vpwr_clk_buf1_branch_0 vpwr_clk_buf1_7 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_8  vpwr_clk_buf1_branch_1 vpwr_clk_buf1_8 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_9  vpwr_clk_buf1_branch_2 vpwr_clk_buf1_9 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_10 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_10 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_11 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_11 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_12 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_12 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_13 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_13 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_14 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_14 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_15 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_15 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_16 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_16 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_17 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_17 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_18 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_18 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_19 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_19 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_20 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_20 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_21 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_21 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_22 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_22 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_23 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_23 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_24 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_24 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_25 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_25 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_26 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_26 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_27 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_27 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_28 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_28 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_29 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_29 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_30 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_30 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_31 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_31 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_32 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_32 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_33 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_33 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_34 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_34 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_35 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_35 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_36 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_36 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_37 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_37 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_38 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_38 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_39 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_39 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_40 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_40 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_41 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_41 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_42 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_42 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_43 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_43 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_44 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_44 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_45 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_45 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_46 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_46 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_47 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_47 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_48 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_48 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_49 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_49 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_50 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_50 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_51 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_51 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_52 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_52 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_53 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_53 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_54 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_54 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_55 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_55 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_56 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_56 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_57 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_57 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_58 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_58 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_59 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_59 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_60 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_60 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_61 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_61 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_62 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_62 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_63 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_63 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_64 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_64 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_65 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_65 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_66 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_66 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_67 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_67 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_68 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_68 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_69 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_69 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_70 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_70 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_71 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_71 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_72 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_72 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_73 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_73 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_74 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_74 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_75 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_75 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_76 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_76 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_77 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_77 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_78 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_78 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_79 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_79 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_80 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_80 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_81 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_81 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_82 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_82 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_83 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_83 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_84 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_84 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_85 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_85 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_86 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_86 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_87 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_87 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_88 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_88 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_89 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_89 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_90 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_90 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_91 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_91 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_92 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_92 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_93 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_93 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_94 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_94 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_95 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_95 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_96 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_96 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_97 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_97 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_98 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_98 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_99 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_99 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_100 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_100 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_101 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_101 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_102 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_102 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_103 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_103 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_104 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_104 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_105 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_105 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_106 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_106 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_107 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_107 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_108 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_108 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_109 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_109 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_110 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_110 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_111 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_111 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_112 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_112 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_113 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_113 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_114 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_114 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_115 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_115 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_116 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_116 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_117 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_117 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_118 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_118 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_119 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_119 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_120 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_120 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_121 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_121 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_122 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_122 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_123 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_123 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_124 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_124 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_125 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_125 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_126 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_126 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_127 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_127 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_128 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_128 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_129 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_129 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_130 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_130 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_131 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_131 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_132 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_132 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_133 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_133 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_134 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_134 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_135 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_135 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_136 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_136 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_137 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_137 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_138 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_138 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_139 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_139 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_140 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_140 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_141 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_141 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_142 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_142 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_143 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_143 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_144 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_144 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_145 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_145 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_146 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_146 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_147 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_147 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_148 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_148 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_149 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_149 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_150 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_150 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_151 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_151 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_152 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_152 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_153 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_153 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_154 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_154 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_155 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_155 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_156 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_156 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_157 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_157 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_158 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_158 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_159 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_159 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_160 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_160 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_161 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_161 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_162 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_162 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_163 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_163 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_164 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_164 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_165 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_165 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_166 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_166 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_167 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_167 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_168 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_168 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_169 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_169 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_170 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_170 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_171 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_171 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_172 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_172 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_173 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_173 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_174 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_174 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_175 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_175 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_176 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_176 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_177 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_177 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_178 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_178 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_179 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_179 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_180 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_180 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_181 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_181 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_182 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_182 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_183 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_183 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_184 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_184 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_185 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_185 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_186 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_186 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_187 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_187 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_188 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_188 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_189 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_189 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_190 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_190 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_191 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_191 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_192 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_192 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_193 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_193 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_194 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_194 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_195 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_195 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_196 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_196 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_197 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_197 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_198 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_198 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_199 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_199 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_200 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_200 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_201 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_201 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_202 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_202 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_203 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_203 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_204 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_204 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_205 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_205 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_206 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_206 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_207 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_207 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_208 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_208 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_209 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_209 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_210 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_210 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_211 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_211 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_212 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_212 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_213 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_213 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_214 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_214 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_215 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_215 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_216 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_216 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_217 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_217 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_218 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_218 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_219 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_219 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_220 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_220 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_221 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_221 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_222 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_222 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_223 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_223 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_224 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_224 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_225 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_225 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_226 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_226 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_227 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_227 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_228 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_228 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_229 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_229 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_230 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_230 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_231 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_231 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_232 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_232 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_233 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_233 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_234 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_234 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_235 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_235 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_236 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_236 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_237 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_237 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_238 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_238 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_239 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_239 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_240 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_240 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_241 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_241 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_242 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_242 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_243 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_243 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_244 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_244 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_245 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_245 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_246 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_246 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_247 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_247 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_248 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_248 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_249 vpwr_clk_buf1_branch_4 vpwr_clk_buf1_249 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_250 vpwr_clk_buf1_branch_5 vpwr_clk_buf1_250 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_251 vpwr_clk_buf1_branch_6 vpwr_clk_buf1_251 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_252 vpwr_clk_buf1_branch_0 vpwr_clk_buf1_252 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_253 vpwr_clk_buf1_branch_1 vpwr_clk_buf1_253 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_254 vpwr_clk_buf1_branch_2 vpwr_clk_buf1_254 ${R_clk_buf1_BUFF}
RP_clk_buf1_LOAD_255 vpwr_clk_buf1_branch_3 vpwr_clk_buf1_255 ${R_clk_buf1_BUFF}
XDC_clk_buf1_0_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_2 VGND VNB vpwr_clk_buf1_2 vpwr_clk_buf1_2 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_2 VGND VNB vpwr_clk_buf1_2 vpwr_clk_buf1_2 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_2 VGND VNB vpwr_clk_buf1_2 vpwr_clk_buf1_2 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_3 VGND VNB vpwr_clk_buf1_3 vpwr_clk_buf1_3 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_3 VGND VNB vpwr_clk_buf1_3 vpwr_clk_buf1_3 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_3 VGND VNB vpwr_clk_buf1_3 vpwr_clk_buf1_3 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_4 VGND VNB vpwr_clk_buf1_4 vpwr_clk_buf1_4 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_4 VGND VNB vpwr_clk_buf1_4 vpwr_clk_buf1_4 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_4 VGND VNB vpwr_clk_buf1_4 vpwr_clk_buf1_4 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_5 VGND VNB vpwr_clk_buf1_5 vpwr_clk_buf1_5 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_5 VGND VNB vpwr_clk_buf1_5 vpwr_clk_buf1_5 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_5 VGND VNB vpwr_clk_buf1_5 vpwr_clk_buf1_5 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_6 VGND VNB vpwr_clk_buf1_6 vpwr_clk_buf1_6 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_6 VGND VNB vpwr_clk_buf1_6 vpwr_clk_buf1_6 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_6 VGND VNB vpwr_clk_buf1_6 vpwr_clk_buf1_6 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_7 VGND VNB vpwr_clk_buf1_7 vpwr_clk_buf1_7 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_7 VGND VNB vpwr_clk_buf1_7 vpwr_clk_buf1_7 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_7 VGND VNB vpwr_clk_buf1_7 vpwr_clk_buf1_7 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_8 VGND VNB vpwr_clk_buf1_8 vpwr_clk_buf1_8 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_8 VGND VNB vpwr_clk_buf1_8 vpwr_clk_buf1_8 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_8 VGND VNB vpwr_clk_buf1_8 vpwr_clk_buf1_8 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_9 VGND VNB vpwr_clk_buf1_9 vpwr_clk_buf1_9 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_9 VGND VNB vpwr_clk_buf1_9 vpwr_clk_buf1_9 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_9 VGND VNB vpwr_clk_buf1_9 vpwr_clk_buf1_9 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_10 VGND VNB vpwr_clk_buf1_10 vpwr_clk_buf1_10 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_10 VGND VNB vpwr_clk_buf1_10 vpwr_clk_buf1_10 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_10 VGND VNB vpwr_clk_buf1_10 vpwr_clk_buf1_10 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_11 VGND VNB vpwr_clk_buf1_11 vpwr_clk_buf1_11 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_11 VGND VNB vpwr_clk_buf1_11 vpwr_clk_buf1_11 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_11 VGND VNB vpwr_clk_buf1_11 vpwr_clk_buf1_11 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_12 VGND VNB vpwr_clk_buf1_12 vpwr_clk_buf1_12 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_12 VGND VNB vpwr_clk_buf1_12 vpwr_clk_buf1_12 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_12 VGND VNB vpwr_clk_buf1_12 vpwr_clk_buf1_12 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_13 VGND VNB vpwr_clk_buf1_13 vpwr_clk_buf1_13 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_13 VGND VNB vpwr_clk_buf1_13 vpwr_clk_buf1_13 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_13 VGND VNB vpwr_clk_buf1_13 vpwr_clk_buf1_13 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_14 VGND VNB vpwr_clk_buf1_14 vpwr_clk_buf1_14 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_14 VGND VNB vpwr_clk_buf1_14 vpwr_clk_buf1_14 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_14 VGND VNB vpwr_clk_buf1_14 vpwr_clk_buf1_14 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_15 VGND VNB vpwr_clk_buf1_15 vpwr_clk_buf1_15 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_15 VGND VNB vpwr_clk_buf1_15 vpwr_clk_buf1_15 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_15 VGND VNB vpwr_clk_buf1_15 vpwr_clk_buf1_15 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_16 VGND VNB vpwr_clk_buf1_16 vpwr_clk_buf1_16 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_16 VGND VNB vpwr_clk_buf1_16 vpwr_clk_buf1_16 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_16 VGND VNB vpwr_clk_buf1_16 vpwr_clk_buf1_16 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_17 VGND VNB vpwr_clk_buf1_17 vpwr_clk_buf1_17 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_17 VGND VNB vpwr_clk_buf1_17 vpwr_clk_buf1_17 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_17 VGND VNB vpwr_clk_buf1_17 vpwr_clk_buf1_17 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_18 VGND VNB vpwr_clk_buf1_18 vpwr_clk_buf1_18 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_18 VGND VNB vpwr_clk_buf1_18 vpwr_clk_buf1_18 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_18 VGND VNB vpwr_clk_buf1_18 vpwr_clk_buf1_18 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_19 VGND VNB vpwr_clk_buf1_19 vpwr_clk_buf1_19 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_19 VGND VNB vpwr_clk_buf1_19 vpwr_clk_buf1_19 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_19 VGND VNB vpwr_clk_buf1_19 vpwr_clk_buf1_19 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_20 VGND VNB vpwr_clk_buf1_20 vpwr_clk_buf1_20 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_20 VGND VNB vpwr_clk_buf1_20 vpwr_clk_buf1_20 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_20 VGND VNB vpwr_clk_buf1_20 vpwr_clk_buf1_20 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_21 VGND VNB vpwr_clk_buf1_21 vpwr_clk_buf1_21 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_21 VGND VNB vpwr_clk_buf1_21 vpwr_clk_buf1_21 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_21 VGND VNB vpwr_clk_buf1_21 vpwr_clk_buf1_21 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_22 VGND VNB vpwr_clk_buf1_22 vpwr_clk_buf1_22 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_22 VGND VNB vpwr_clk_buf1_22 vpwr_clk_buf1_22 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_22 VGND VNB vpwr_clk_buf1_22 vpwr_clk_buf1_22 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_23 VGND VNB vpwr_clk_buf1_23 vpwr_clk_buf1_23 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_23 VGND VNB vpwr_clk_buf1_23 vpwr_clk_buf1_23 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_23 VGND VNB vpwr_clk_buf1_23 vpwr_clk_buf1_23 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_24 VGND VNB vpwr_clk_buf1_24 vpwr_clk_buf1_24 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_24 VGND VNB vpwr_clk_buf1_24 vpwr_clk_buf1_24 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_24 VGND VNB vpwr_clk_buf1_24 vpwr_clk_buf1_24 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_25 VGND VNB vpwr_clk_buf1_25 vpwr_clk_buf1_25 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_25 VGND VNB vpwr_clk_buf1_25 vpwr_clk_buf1_25 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_25 VGND VNB vpwr_clk_buf1_25 vpwr_clk_buf1_25 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_26 VGND VNB vpwr_clk_buf1_26 vpwr_clk_buf1_26 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_26 VGND VNB vpwr_clk_buf1_26 vpwr_clk_buf1_26 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_26 VGND VNB vpwr_clk_buf1_26 vpwr_clk_buf1_26 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_27 VGND VNB vpwr_clk_buf1_27 vpwr_clk_buf1_27 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_27 VGND VNB vpwr_clk_buf1_27 vpwr_clk_buf1_27 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_27 VGND VNB vpwr_clk_buf1_27 vpwr_clk_buf1_27 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_28 VGND VNB vpwr_clk_buf1_28 vpwr_clk_buf1_28 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_28 VGND VNB vpwr_clk_buf1_28 vpwr_clk_buf1_28 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_28 VGND VNB vpwr_clk_buf1_28 vpwr_clk_buf1_28 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_29 VGND VNB vpwr_clk_buf1_29 vpwr_clk_buf1_29 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_29 VGND VNB vpwr_clk_buf1_29 vpwr_clk_buf1_29 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_29 VGND VNB vpwr_clk_buf1_29 vpwr_clk_buf1_29 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_30 VGND VNB vpwr_clk_buf1_30 vpwr_clk_buf1_30 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_30 VGND VNB vpwr_clk_buf1_30 vpwr_clk_buf1_30 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_30 VGND VNB vpwr_clk_buf1_30 vpwr_clk_buf1_30 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_31 VGND VNB vpwr_clk_buf1_31 vpwr_clk_buf1_31 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_31 VGND VNB vpwr_clk_buf1_31 vpwr_clk_buf1_31 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_31 VGND VNB vpwr_clk_buf1_31 vpwr_clk_buf1_31 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_32 VGND VNB vpwr_clk_buf1_32 vpwr_clk_buf1_32 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_32 VGND VNB vpwr_clk_buf1_32 vpwr_clk_buf1_32 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_32 VGND VNB vpwr_clk_buf1_32 vpwr_clk_buf1_32 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_33 VGND VNB vpwr_clk_buf1_33 vpwr_clk_buf1_33 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_33 VGND VNB vpwr_clk_buf1_33 vpwr_clk_buf1_33 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_33 VGND VNB vpwr_clk_buf1_33 vpwr_clk_buf1_33 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_34 VGND VNB vpwr_clk_buf1_34 vpwr_clk_buf1_34 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_34 VGND VNB vpwr_clk_buf1_34 vpwr_clk_buf1_34 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_34 VGND VNB vpwr_clk_buf1_34 vpwr_clk_buf1_34 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_35 VGND VNB vpwr_clk_buf1_35 vpwr_clk_buf1_35 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_35 VGND VNB vpwr_clk_buf1_35 vpwr_clk_buf1_35 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_35 VGND VNB vpwr_clk_buf1_35 vpwr_clk_buf1_35 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_36 VGND VNB vpwr_clk_buf1_36 vpwr_clk_buf1_36 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_36 VGND VNB vpwr_clk_buf1_36 vpwr_clk_buf1_36 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_36 VGND VNB vpwr_clk_buf1_36 vpwr_clk_buf1_36 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_37 VGND VNB vpwr_clk_buf1_37 vpwr_clk_buf1_37 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_37 VGND VNB vpwr_clk_buf1_37 vpwr_clk_buf1_37 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_37 VGND VNB vpwr_clk_buf1_37 vpwr_clk_buf1_37 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_38 VGND VNB vpwr_clk_buf1_38 vpwr_clk_buf1_38 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_38 VGND VNB vpwr_clk_buf1_38 vpwr_clk_buf1_38 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_38 VGND VNB vpwr_clk_buf1_38 vpwr_clk_buf1_38 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_39 VGND VNB vpwr_clk_buf1_39 vpwr_clk_buf1_39 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_39 VGND VNB vpwr_clk_buf1_39 vpwr_clk_buf1_39 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_39 VGND VNB vpwr_clk_buf1_39 vpwr_clk_buf1_39 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_40 VGND VNB vpwr_clk_buf1_40 vpwr_clk_buf1_40 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_40 VGND VNB vpwr_clk_buf1_40 vpwr_clk_buf1_40 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_40 VGND VNB vpwr_clk_buf1_40 vpwr_clk_buf1_40 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_41 VGND VNB vpwr_clk_buf1_41 vpwr_clk_buf1_41 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_41 VGND VNB vpwr_clk_buf1_41 vpwr_clk_buf1_41 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_41 VGND VNB vpwr_clk_buf1_41 vpwr_clk_buf1_41 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_42 VGND VNB vpwr_clk_buf1_42 vpwr_clk_buf1_42 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_42 VGND VNB vpwr_clk_buf1_42 vpwr_clk_buf1_42 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_42 VGND VNB vpwr_clk_buf1_42 vpwr_clk_buf1_42 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_43 VGND VNB vpwr_clk_buf1_43 vpwr_clk_buf1_43 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_43 VGND VNB vpwr_clk_buf1_43 vpwr_clk_buf1_43 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_43 VGND VNB vpwr_clk_buf1_43 vpwr_clk_buf1_43 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_44 VGND VNB vpwr_clk_buf1_44 vpwr_clk_buf1_44 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_44 VGND VNB vpwr_clk_buf1_44 vpwr_clk_buf1_44 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_44 VGND VNB vpwr_clk_buf1_44 vpwr_clk_buf1_44 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_45 VGND VNB vpwr_clk_buf1_45 vpwr_clk_buf1_45 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_45 VGND VNB vpwr_clk_buf1_45 vpwr_clk_buf1_45 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_45 VGND VNB vpwr_clk_buf1_45 vpwr_clk_buf1_45 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_46 VGND VNB vpwr_clk_buf1_46 vpwr_clk_buf1_46 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_46 VGND VNB vpwr_clk_buf1_46 vpwr_clk_buf1_46 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_46 VGND VNB vpwr_clk_buf1_46 vpwr_clk_buf1_46 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_47 VGND VNB vpwr_clk_buf1_47 vpwr_clk_buf1_47 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_47 VGND VNB vpwr_clk_buf1_47 vpwr_clk_buf1_47 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_47 VGND VNB vpwr_clk_buf1_47 vpwr_clk_buf1_47 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_48 VGND VNB vpwr_clk_buf1_48 vpwr_clk_buf1_48 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_48 VGND VNB vpwr_clk_buf1_48 vpwr_clk_buf1_48 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_48 VGND VNB vpwr_clk_buf1_48 vpwr_clk_buf1_48 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_49 VGND VNB vpwr_clk_buf1_49 vpwr_clk_buf1_49 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_49 VGND VNB vpwr_clk_buf1_49 vpwr_clk_buf1_49 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_49 VGND VNB vpwr_clk_buf1_49 vpwr_clk_buf1_49 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_50 VGND VNB vpwr_clk_buf1_50 vpwr_clk_buf1_50 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_50 VGND VNB vpwr_clk_buf1_50 vpwr_clk_buf1_50 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_50 VGND VNB vpwr_clk_buf1_50 vpwr_clk_buf1_50 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_51 VGND VNB vpwr_clk_buf1_51 vpwr_clk_buf1_51 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_51 VGND VNB vpwr_clk_buf1_51 vpwr_clk_buf1_51 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_51 VGND VNB vpwr_clk_buf1_51 vpwr_clk_buf1_51 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_52 VGND VNB vpwr_clk_buf1_52 vpwr_clk_buf1_52 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_52 VGND VNB vpwr_clk_buf1_52 vpwr_clk_buf1_52 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_52 VGND VNB vpwr_clk_buf1_52 vpwr_clk_buf1_52 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_53 VGND VNB vpwr_clk_buf1_53 vpwr_clk_buf1_53 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_53 VGND VNB vpwr_clk_buf1_53 vpwr_clk_buf1_53 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_53 VGND VNB vpwr_clk_buf1_53 vpwr_clk_buf1_53 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_54 VGND VNB vpwr_clk_buf1_54 vpwr_clk_buf1_54 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_54 VGND VNB vpwr_clk_buf1_54 vpwr_clk_buf1_54 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_54 VGND VNB vpwr_clk_buf1_54 vpwr_clk_buf1_54 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_55 VGND VNB vpwr_clk_buf1_55 vpwr_clk_buf1_55 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_55 VGND VNB vpwr_clk_buf1_55 vpwr_clk_buf1_55 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_55 VGND VNB vpwr_clk_buf1_55 vpwr_clk_buf1_55 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_56 VGND VNB vpwr_clk_buf1_56 vpwr_clk_buf1_56 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_56 VGND VNB vpwr_clk_buf1_56 vpwr_clk_buf1_56 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_56 VGND VNB vpwr_clk_buf1_56 vpwr_clk_buf1_56 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_57 VGND VNB vpwr_clk_buf1_57 vpwr_clk_buf1_57 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_57 VGND VNB vpwr_clk_buf1_57 vpwr_clk_buf1_57 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_57 VGND VNB vpwr_clk_buf1_57 vpwr_clk_buf1_57 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_58 VGND VNB vpwr_clk_buf1_58 vpwr_clk_buf1_58 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_58 VGND VNB vpwr_clk_buf1_58 vpwr_clk_buf1_58 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_58 VGND VNB vpwr_clk_buf1_58 vpwr_clk_buf1_58 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_59 VGND VNB vpwr_clk_buf1_59 vpwr_clk_buf1_59 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_59 VGND VNB vpwr_clk_buf1_59 vpwr_clk_buf1_59 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_59 VGND VNB vpwr_clk_buf1_59 vpwr_clk_buf1_59 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_60 VGND VNB vpwr_clk_buf1_60 vpwr_clk_buf1_60 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_60 VGND VNB vpwr_clk_buf1_60 vpwr_clk_buf1_60 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_60 VGND VNB vpwr_clk_buf1_60 vpwr_clk_buf1_60 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_61 VGND VNB vpwr_clk_buf1_61 vpwr_clk_buf1_61 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_61 VGND VNB vpwr_clk_buf1_61 vpwr_clk_buf1_61 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_61 VGND VNB vpwr_clk_buf1_61 vpwr_clk_buf1_61 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_62 VGND VNB vpwr_clk_buf1_62 vpwr_clk_buf1_62 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_62 VGND VNB vpwr_clk_buf1_62 vpwr_clk_buf1_62 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_62 VGND VNB vpwr_clk_buf1_62 vpwr_clk_buf1_62 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_63 VGND VNB vpwr_clk_buf1_63 vpwr_clk_buf1_63 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_63 VGND VNB vpwr_clk_buf1_63 vpwr_clk_buf1_63 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_63 VGND VNB vpwr_clk_buf1_63 vpwr_clk_buf1_63 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_64 VGND VNB vpwr_clk_buf1_64 vpwr_clk_buf1_64 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_64 VGND VNB vpwr_clk_buf1_64 vpwr_clk_buf1_64 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_64 VGND VNB vpwr_clk_buf1_64 vpwr_clk_buf1_64 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_65 VGND VNB vpwr_clk_buf1_65 vpwr_clk_buf1_65 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_65 VGND VNB vpwr_clk_buf1_65 vpwr_clk_buf1_65 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_65 VGND VNB vpwr_clk_buf1_65 vpwr_clk_buf1_65 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_66 VGND VNB vpwr_clk_buf1_66 vpwr_clk_buf1_66 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_66 VGND VNB vpwr_clk_buf1_66 vpwr_clk_buf1_66 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_66 VGND VNB vpwr_clk_buf1_66 vpwr_clk_buf1_66 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_67 VGND VNB vpwr_clk_buf1_67 vpwr_clk_buf1_67 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_67 VGND VNB vpwr_clk_buf1_67 vpwr_clk_buf1_67 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_67 VGND VNB vpwr_clk_buf1_67 vpwr_clk_buf1_67 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_68 VGND VNB vpwr_clk_buf1_68 vpwr_clk_buf1_68 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_68 VGND VNB vpwr_clk_buf1_68 vpwr_clk_buf1_68 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_68 VGND VNB vpwr_clk_buf1_68 vpwr_clk_buf1_68 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_69 VGND VNB vpwr_clk_buf1_69 vpwr_clk_buf1_69 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_69 VGND VNB vpwr_clk_buf1_69 vpwr_clk_buf1_69 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_69 VGND VNB vpwr_clk_buf1_69 vpwr_clk_buf1_69 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_70 VGND VNB vpwr_clk_buf1_70 vpwr_clk_buf1_70 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_70 VGND VNB vpwr_clk_buf1_70 vpwr_clk_buf1_70 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_70 VGND VNB vpwr_clk_buf1_70 vpwr_clk_buf1_70 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_71 VGND VNB vpwr_clk_buf1_71 vpwr_clk_buf1_71 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_71 VGND VNB vpwr_clk_buf1_71 vpwr_clk_buf1_71 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_71 VGND VNB vpwr_clk_buf1_71 vpwr_clk_buf1_71 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_72 VGND VNB vpwr_clk_buf1_72 vpwr_clk_buf1_72 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_72 VGND VNB vpwr_clk_buf1_72 vpwr_clk_buf1_72 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_72 VGND VNB vpwr_clk_buf1_72 vpwr_clk_buf1_72 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_73 VGND VNB vpwr_clk_buf1_73 vpwr_clk_buf1_73 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_73 VGND VNB vpwr_clk_buf1_73 vpwr_clk_buf1_73 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_73 VGND VNB vpwr_clk_buf1_73 vpwr_clk_buf1_73 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_74 VGND VNB vpwr_clk_buf1_74 vpwr_clk_buf1_74 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_74 VGND VNB vpwr_clk_buf1_74 vpwr_clk_buf1_74 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_74 VGND VNB vpwr_clk_buf1_74 vpwr_clk_buf1_74 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_75 VGND VNB vpwr_clk_buf1_75 vpwr_clk_buf1_75 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_75 VGND VNB vpwr_clk_buf1_75 vpwr_clk_buf1_75 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_75 VGND VNB vpwr_clk_buf1_75 vpwr_clk_buf1_75 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_76 VGND VNB vpwr_clk_buf1_76 vpwr_clk_buf1_76 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_76 VGND VNB vpwr_clk_buf1_76 vpwr_clk_buf1_76 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_76 VGND VNB vpwr_clk_buf1_76 vpwr_clk_buf1_76 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_77 VGND VNB vpwr_clk_buf1_77 vpwr_clk_buf1_77 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_77 VGND VNB vpwr_clk_buf1_77 vpwr_clk_buf1_77 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_77 VGND VNB vpwr_clk_buf1_77 vpwr_clk_buf1_77 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_78 VGND VNB vpwr_clk_buf1_78 vpwr_clk_buf1_78 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_78 VGND VNB vpwr_clk_buf1_78 vpwr_clk_buf1_78 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_78 VGND VNB vpwr_clk_buf1_78 vpwr_clk_buf1_78 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_79 VGND VNB vpwr_clk_buf1_79 vpwr_clk_buf1_79 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_79 VGND VNB vpwr_clk_buf1_79 vpwr_clk_buf1_79 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_79 VGND VNB vpwr_clk_buf1_79 vpwr_clk_buf1_79 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_80 VGND VNB vpwr_clk_buf1_80 vpwr_clk_buf1_80 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_80 VGND VNB vpwr_clk_buf1_80 vpwr_clk_buf1_80 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_80 VGND VNB vpwr_clk_buf1_80 vpwr_clk_buf1_80 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_81 VGND VNB vpwr_clk_buf1_81 vpwr_clk_buf1_81 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_81 VGND VNB vpwr_clk_buf1_81 vpwr_clk_buf1_81 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_81 VGND VNB vpwr_clk_buf1_81 vpwr_clk_buf1_81 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_82 VGND VNB vpwr_clk_buf1_82 vpwr_clk_buf1_82 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_82 VGND VNB vpwr_clk_buf1_82 vpwr_clk_buf1_82 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_82 VGND VNB vpwr_clk_buf1_82 vpwr_clk_buf1_82 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_83 VGND VNB vpwr_clk_buf1_83 vpwr_clk_buf1_83 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_83 VGND VNB vpwr_clk_buf1_83 vpwr_clk_buf1_83 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_83 VGND VNB vpwr_clk_buf1_83 vpwr_clk_buf1_83 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_84 VGND VNB vpwr_clk_buf1_84 vpwr_clk_buf1_84 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_84 VGND VNB vpwr_clk_buf1_84 vpwr_clk_buf1_84 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_84 VGND VNB vpwr_clk_buf1_84 vpwr_clk_buf1_84 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_85 VGND VNB vpwr_clk_buf1_85 vpwr_clk_buf1_85 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_85 VGND VNB vpwr_clk_buf1_85 vpwr_clk_buf1_85 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_85 VGND VNB vpwr_clk_buf1_85 vpwr_clk_buf1_85 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_86 VGND VNB vpwr_clk_buf1_86 vpwr_clk_buf1_86 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_86 VGND VNB vpwr_clk_buf1_86 vpwr_clk_buf1_86 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_86 VGND VNB vpwr_clk_buf1_86 vpwr_clk_buf1_86 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_87 VGND VNB vpwr_clk_buf1_87 vpwr_clk_buf1_87 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_87 VGND VNB vpwr_clk_buf1_87 vpwr_clk_buf1_87 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_87 VGND VNB vpwr_clk_buf1_87 vpwr_clk_buf1_87 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_88 VGND VNB vpwr_clk_buf1_88 vpwr_clk_buf1_88 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_88 VGND VNB vpwr_clk_buf1_88 vpwr_clk_buf1_88 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_88 VGND VNB vpwr_clk_buf1_88 vpwr_clk_buf1_88 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_89 VGND VNB vpwr_clk_buf1_89 vpwr_clk_buf1_89 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_89 VGND VNB vpwr_clk_buf1_89 vpwr_clk_buf1_89 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_89 VGND VNB vpwr_clk_buf1_89 vpwr_clk_buf1_89 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_90 VGND VNB vpwr_clk_buf1_90 vpwr_clk_buf1_90 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_90 VGND VNB vpwr_clk_buf1_90 vpwr_clk_buf1_90 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_90 VGND VNB vpwr_clk_buf1_90 vpwr_clk_buf1_90 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_91 VGND VNB vpwr_clk_buf1_91 vpwr_clk_buf1_91 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_91 VGND VNB vpwr_clk_buf1_91 vpwr_clk_buf1_91 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_91 VGND VNB vpwr_clk_buf1_91 vpwr_clk_buf1_91 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_92 VGND VNB vpwr_clk_buf1_92 vpwr_clk_buf1_92 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_92 VGND VNB vpwr_clk_buf1_92 vpwr_clk_buf1_92 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_92 VGND VNB vpwr_clk_buf1_92 vpwr_clk_buf1_92 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_93 VGND VNB vpwr_clk_buf1_93 vpwr_clk_buf1_93 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_93 VGND VNB vpwr_clk_buf1_93 vpwr_clk_buf1_93 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_93 VGND VNB vpwr_clk_buf1_93 vpwr_clk_buf1_93 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_94 VGND VNB vpwr_clk_buf1_94 vpwr_clk_buf1_94 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_94 VGND VNB vpwr_clk_buf1_94 vpwr_clk_buf1_94 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_94 VGND VNB vpwr_clk_buf1_94 vpwr_clk_buf1_94 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_95 VGND VNB vpwr_clk_buf1_95 vpwr_clk_buf1_95 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_95 VGND VNB vpwr_clk_buf1_95 vpwr_clk_buf1_95 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_95 VGND VNB vpwr_clk_buf1_95 vpwr_clk_buf1_95 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_96 VGND VNB vpwr_clk_buf1_96 vpwr_clk_buf1_96 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_96 VGND VNB vpwr_clk_buf1_96 vpwr_clk_buf1_96 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_96 VGND VNB vpwr_clk_buf1_96 vpwr_clk_buf1_96 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_97 VGND VNB vpwr_clk_buf1_97 vpwr_clk_buf1_97 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_97 VGND VNB vpwr_clk_buf1_97 vpwr_clk_buf1_97 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_97 VGND VNB vpwr_clk_buf1_97 vpwr_clk_buf1_97 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_98 VGND VNB vpwr_clk_buf1_98 vpwr_clk_buf1_98 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_98 VGND VNB vpwr_clk_buf1_98 vpwr_clk_buf1_98 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_98 VGND VNB vpwr_clk_buf1_98 vpwr_clk_buf1_98 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_99 VGND VNB vpwr_clk_buf1_99 vpwr_clk_buf1_99 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_99 VGND VNB vpwr_clk_buf1_99 vpwr_clk_buf1_99 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_99 VGND VNB vpwr_clk_buf1_99 vpwr_clk_buf1_99 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_100 VGND VNB vpwr_clk_buf1_100 vpwr_clk_buf1_100 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_100 VGND VNB vpwr_clk_buf1_100 vpwr_clk_buf1_100 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_100 VGND VNB vpwr_clk_buf1_100 vpwr_clk_buf1_100 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_101 VGND VNB vpwr_clk_buf1_101 vpwr_clk_buf1_101 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_101 VGND VNB vpwr_clk_buf1_101 vpwr_clk_buf1_101 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_101 VGND VNB vpwr_clk_buf1_101 vpwr_clk_buf1_101 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_102 VGND VNB vpwr_clk_buf1_102 vpwr_clk_buf1_102 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_102 VGND VNB vpwr_clk_buf1_102 vpwr_clk_buf1_102 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_102 VGND VNB vpwr_clk_buf1_102 vpwr_clk_buf1_102 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_103 VGND VNB vpwr_clk_buf1_103 vpwr_clk_buf1_103 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_103 VGND VNB vpwr_clk_buf1_103 vpwr_clk_buf1_103 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_103 VGND VNB vpwr_clk_buf1_103 vpwr_clk_buf1_103 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_104 VGND VNB vpwr_clk_buf1_104 vpwr_clk_buf1_104 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_104 VGND VNB vpwr_clk_buf1_104 vpwr_clk_buf1_104 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_104 VGND VNB vpwr_clk_buf1_104 vpwr_clk_buf1_104 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_105 VGND VNB vpwr_clk_buf1_105 vpwr_clk_buf1_105 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_105 VGND VNB vpwr_clk_buf1_105 vpwr_clk_buf1_105 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_105 VGND VNB vpwr_clk_buf1_105 vpwr_clk_buf1_105 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_106 VGND VNB vpwr_clk_buf1_106 vpwr_clk_buf1_106 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_106 VGND VNB vpwr_clk_buf1_106 vpwr_clk_buf1_106 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_106 VGND VNB vpwr_clk_buf1_106 vpwr_clk_buf1_106 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_107 VGND VNB vpwr_clk_buf1_107 vpwr_clk_buf1_107 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_107 VGND VNB vpwr_clk_buf1_107 vpwr_clk_buf1_107 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_107 VGND VNB vpwr_clk_buf1_107 vpwr_clk_buf1_107 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_108 VGND VNB vpwr_clk_buf1_108 vpwr_clk_buf1_108 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_108 VGND VNB vpwr_clk_buf1_108 vpwr_clk_buf1_108 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_108 VGND VNB vpwr_clk_buf1_108 vpwr_clk_buf1_108 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_109 VGND VNB vpwr_clk_buf1_109 vpwr_clk_buf1_109 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_109 VGND VNB vpwr_clk_buf1_109 vpwr_clk_buf1_109 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_109 VGND VNB vpwr_clk_buf1_109 vpwr_clk_buf1_109 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_110 VGND VNB vpwr_clk_buf1_110 vpwr_clk_buf1_110 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_110 VGND VNB vpwr_clk_buf1_110 vpwr_clk_buf1_110 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_110 VGND VNB vpwr_clk_buf1_110 vpwr_clk_buf1_110 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_111 VGND VNB vpwr_clk_buf1_111 vpwr_clk_buf1_111 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_111 VGND VNB vpwr_clk_buf1_111 vpwr_clk_buf1_111 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_111 VGND VNB vpwr_clk_buf1_111 vpwr_clk_buf1_111 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_112 VGND VNB vpwr_clk_buf1_112 vpwr_clk_buf1_112 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_112 VGND VNB vpwr_clk_buf1_112 vpwr_clk_buf1_112 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_112 VGND VNB vpwr_clk_buf1_112 vpwr_clk_buf1_112 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_113 VGND VNB vpwr_clk_buf1_113 vpwr_clk_buf1_113 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_113 VGND VNB vpwr_clk_buf1_113 vpwr_clk_buf1_113 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_113 VGND VNB vpwr_clk_buf1_113 vpwr_clk_buf1_113 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_114 VGND VNB vpwr_clk_buf1_114 vpwr_clk_buf1_114 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_114 VGND VNB vpwr_clk_buf1_114 vpwr_clk_buf1_114 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_114 VGND VNB vpwr_clk_buf1_114 vpwr_clk_buf1_114 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_115 VGND VNB vpwr_clk_buf1_115 vpwr_clk_buf1_115 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_115 VGND VNB vpwr_clk_buf1_115 vpwr_clk_buf1_115 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_115 VGND VNB vpwr_clk_buf1_115 vpwr_clk_buf1_115 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_116 VGND VNB vpwr_clk_buf1_116 vpwr_clk_buf1_116 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_116 VGND VNB vpwr_clk_buf1_116 vpwr_clk_buf1_116 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_116 VGND VNB vpwr_clk_buf1_116 vpwr_clk_buf1_116 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_117 VGND VNB vpwr_clk_buf1_117 vpwr_clk_buf1_117 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_117 VGND VNB vpwr_clk_buf1_117 vpwr_clk_buf1_117 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_117 VGND VNB vpwr_clk_buf1_117 vpwr_clk_buf1_117 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_118 VGND VNB vpwr_clk_buf1_118 vpwr_clk_buf1_118 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_118 VGND VNB vpwr_clk_buf1_118 vpwr_clk_buf1_118 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_118 VGND VNB vpwr_clk_buf1_118 vpwr_clk_buf1_118 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_119 VGND VNB vpwr_clk_buf1_119 vpwr_clk_buf1_119 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_119 VGND VNB vpwr_clk_buf1_119 vpwr_clk_buf1_119 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_119 VGND VNB vpwr_clk_buf1_119 vpwr_clk_buf1_119 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_120 VGND VNB vpwr_clk_buf1_120 vpwr_clk_buf1_120 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_120 VGND VNB vpwr_clk_buf1_120 vpwr_clk_buf1_120 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_120 VGND VNB vpwr_clk_buf1_120 vpwr_clk_buf1_120 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_121 VGND VNB vpwr_clk_buf1_121 vpwr_clk_buf1_121 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_121 VGND VNB vpwr_clk_buf1_121 vpwr_clk_buf1_121 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_121 VGND VNB vpwr_clk_buf1_121 vpwr_clk_buf1_121 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_122 VGND VNB vpwr_clk_buf1_122 vpwr_clk_buf1_122 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_122 VGND VNB vpwr_clk_buf1_122 vpwr_clk_buf1_122 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_122 VGND VNB vpwr_clk_buf1_122 vpwr_clk_buf1_122 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_123 VGND VNB vpwr_clk_buf1_123 vpwr_clk_buf1_123 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_123 VGND VNB vpwr_clk_buf1_123 vpwr_clk_buf1_123 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_123 VGND VNB vpwr_clk_buf1_123 vpwr_clk_buf1_123 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_124 VGND VNB vpwr_clk_buf1_124 vpwr_clk_buf1_124 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_124 VGND VNB vpwr_clk_buf1_124 vpwr_clk_buf1_124 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_124 VGND VNB vpwr_clk_buf1_124 vpwr_clk_buf1_124 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_125 VGND VNB vpwr_clk_buf1_125 vpwr_clk_buf1_125 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_125 VGND VNB vpwr_clk_buf1_125 vpwr_clk_buf1_125 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_125 VGND VNB vpwr_clk_buf1_125 vpwr_clk_buf1_125 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_126 VGND VNB vpwr_clk_buf1_126 vpwr_clk_buf1_126 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_126 VGND VNB vpwr_clk_buf1_126 vpwr_clk_buf1_126 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_126 VGND VNB vpwr_clk_buf1_126 vpwr_clk_buf1_126 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_127 VGND VNB vpwr_clk_buf1_127 vpwr_clk_buf1_127 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_127 VGND VNB vpwr_clk_buf1_127 vpwr_clk_buf1_127 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_127 VGND VNB vpwr_clk_buf1_127 vpwr_clk_buf1_127 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_128 VGND VNB vpwr_clk_buf1_128 vpwr_clk_buf1_128 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_128 VGND VNB vpwr_clk_buf1_128 vpwr_clk_buf1_128 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_128 VGND VNB vpwr_clk_buf1_128 vpwr_clk_buf1_128 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_129 VGND VNB vpwr_clk_buf1_129 vpwr_clk_buf1_129 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_129 VGND VNB vpwr_clk_buf1_129 vpwr_clk_buf1_129 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_129 VGND VNB vpwr_clk_buf1_129 vpwr_clk_buf1_129 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_130 VGND VNB vpwr_clk_buf1_130 vpwr_clk_buf1_130 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_130 VGND VNB vpwr_clk_buf1_130 vpwr_clk_buf1_130 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_130 VGND VNB vpwr_clk_buf1_130 vpwr_clk_buf1_130 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_131 VGND VNB vpwr_clk_buf1_131 vpwr_clk_buf1_131 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_131 VGND VNB vpwr_clk_buf1_131 vpwr_clk_buf1_131 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_131 VGND VNB vpwr_clk_buf1_131 vpwr_clk_buf1_131 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_132 VGND VNB vpwr_clk_buf1_132 vpwr_clk_buf1_132 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_132 VGND VNB vpwr_clk_buf1_132 vpwr_clk_buf1_132 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_132 VGND VNB vpwr_clk_buf1_132 vpwr_clk_buf1_132 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_133 VGND VNB vpwr_clk_buf1_133 vpwr_clk_buf1_133 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_133 VGND VNB vpwr_clk_buf1_133 vpwr_clk_buf1_133 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_133 VGND VNB vpwr_clk_buf1_133 vpwr_clk_buf1_133 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_134 VGND VNB vpwr_clk_buf1_134 vpwr_clk_buf1_134 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_134 VGND VNB vpwr_clk_buf1_134 vpwr_clk_buf1_134 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_134 VGND VNB vpwr_clk_buf1_134 vpwr_clk_buf1_134 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_135 VGND VNB vpwr_clk_buf1_135 vpwr_clk_buf1_135 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_135 VGND VNB vpwr_clk_buf1_135 vpwr_clk_buf1_135 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_135 VGND VNB vpwr_clk_buf1_135 vpwr_clk_buf1_135 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_136 VGND VNB vpwr_clk_buf1_136 vpwr_clk_buf1_136 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_136 VGND VNB vpwr_clk_buf1_136 vpwr_clk_buf1_136 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_136 VGND VNB vpwr_clk_buf1_136 vpwr_clk_buf1_136 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_137 VGND VNB vpwr_clk_buf1_137 vpwr_clk_buf1_137 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_137 VGND VNB vpwr_clk_buf1_137 vpwr_clk_buf1_137 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_137 VGND VNB vpwr_clk_buf1_137 vpwr_clk_buf1_137 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_138 VGND VNB vpwr_clk_buf1_138 vpwr_clk_buf1_138 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_138 VGND VNB vpwr_clk_buf1_138 vpwr_clk_buf1_138 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_138 VGND VNB vpwr_clk_buf1_138 vpwr_clk_buf1_138 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_139 VGND VNB vpwr_clk_buf1_139 vpwr_clk_buf1_139 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_139 VGND VNB vpwr_clk_buf1_139 vpwr_clk_buf1_139 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_139 VGND VNB vpwr_clk_buf1_139 vpwr_clk_buf1_139 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_140 VGND VNB vpwr_clk_buf1_140 vpwr_clk_buf1_140 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_140 VGND VNB vpwr_clk_buf1_140 vpwr_clk_buf1_140 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_140 VGND VNB vpwr_clk_buf1_140 vpwr_clk_buf1_140 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_141 VGND VNB vpwr_clk_buf1_141 vpwr_clk_buf1_141 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_141 VGND VNB vpwr_clk_buf1_141 vpwr_clk_buf1_141 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_141 VGND VNB vpwr_clk_buf1_141 vpwr_clk_buf1_141 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_142 VGND VNB vpwr_clk_buf1_142 vpwr_clk_buf1_142 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_142 VGND VNB vpwr_clk_buf1_142 vpwr_clk_buf1_142 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_142 VGND VNB vpwr_clk_buf1_142 vpwr_clk_buf1_142 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_143 VGND VNB vpwr_clk_buf1_143 vpwr_clk_buf1_143 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_143 VGND VNB vpwr_clk_buf1_143 vpwr_clk_buf1_143 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_143 VGND VNB vpwr_clk_buf1_143 vpwr_clk_buf1_143 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_144 VGND VNB vpwr_clk_buf1_144 vpwr_clk_buf1_144 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_144 VGND VNB vpwr_clk_buf1_144 vpwr_clk_buf1_144 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_144 VGND VNB vpwr_clk_buf1_144 vpwr_clk_buf1_144 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_145 VGND VNB vpwr_clk_buf1_145 vpwr_clk_buf1_145 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_145 VGND VNB vpwr_clk_buf1_145 vpwr_clk_buf1_145 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_145 VGND VNB vpwr_clk_buf1_145 vpwr_clk_buf1_145 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_146 VGND VNB vpwr_clk_buf1_146 vpwr_clk_buf1_146 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_146 VGND VNB vpwr_clk_buf1_146 vpwr_clk_buf1_146 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_146 VGND VNB vpwr_clk_buf1_146 vpwr_clk_buf1_146 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_147 VGND VNB vpwr_clk_buf1_147 vpwr_clk_buf1_147 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_147 VGND VNB vpwr_clk_buf1_147 vpwr_clk_buf1_147 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_147 VGND VNB vpwr_clk_buf1_147 vpwr_clk_buf1_147 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_148 VGND VNB vpwr_clk_buf1_148 vpwr_clk_buf1_148 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_148 VGND VNB vpwr_clk_buf1_148 vpwr_clk_buf1_148 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_148 VGND VNB vpwr_clk_buf1_148 vpwr_clk_buf1_148 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_149 VGND VNB vpwr_clk_buf1_149 vpwr_clk_buf1_149 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_149 VGND VNB vpwr_clk_buf1_149 vpwr_clk_buf1_149 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_149 VGND VNB vpwr_clk_buf1_149 vpwr_clk_buf1_149 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_150 VGND VNB vpwr_clk_buf1_150 vpwr_clk_buf1_150 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_150 VGND VNB vpwr_clk_buf1_150 vpwr_clk_buf1_150 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_150 VGND VNB vpwr_clk_buf1_150 vpwr_clk_buf1_150 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_151 VGND VNB vpwr_clk_buf1_151 vpwr_clk_buf1_151 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_151 VGND VNB vpwr_clk_buf1_151 vpwr_clk_buf1_151 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_151 VGND VNB vpwr_clk_buf1_151 vpwr_clk_buf1_151 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_152 VGND VNB vpwr_clk_buf1_152 vpwr_clk_buf1_152 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_152 VGND VNB vpwr_clk_buf1_152 vpwr_clk_buf1_152 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_152 VGND VNB vpwr_clk_buf1_152 vpwr_clk_buf1_152 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_153 VGND VNB vpwr_clk_buf1_153 vpwr_clk_buf1_153 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_153 VGND VNB vpwr_clk_buf1_153 vpwr_clk_buf1_153 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_153 VGND VNB vpwr_clk_buf1_153 vpwr_clk_buf1_153 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_154 VGND VNB vpwr_clk_buf1_154 vpwr_clk_buf1_154 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_154 VGND VNB vpwr_clk_buf1_154 vpwr_clk_buf1_154 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_154 VGND VNB vpwr_clk_buf1_154 vpwr_clk_buf1_154 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_155 VGND VNB vpwr_clk_buf1_155 vpwr_clk_buf1_155 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_155 VGND VNB vpwr_clk_buf1_155 vpwr_clk_buf1_155 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_155 VGND VNB vpwr_clk_buf1_155 vpwr_clk_buf1_155 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_156 VGND VNB vpwr_clk_buf1_156 vpwr_clk_buf1_156 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_156 VGND VNB vpwr_clk_buf1_156 vpwr_clk_buf1_156 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_156 VGND VNB vpwr_clk_buf1_156 vpwr_clk_buf1_156 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_157 VGND VNB vpwr_clk_buf1_157 vpwr_clk_buf1_157 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_157 VGND VNB vpwr_clk_buf1_157 vpwr_clk_buf1_157 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_157 VGND VNB vpwr_clk_buf1_157 vpwr_clk_buf1_157 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_158 VGND VNB vpwr_clk_buf1_158 vpwr_clk_buf1_158 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_158 VGND VNB vpwr_clk_buf1_158 vpwr_clk_buf1_158 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_158 VGND VNB vpwr_clk_buf1_158 vpwr_clk_buf1_158 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_159 VGND VNB vpwr_clk_buf1_159 vpwr_clk_buf1_159 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_159 VGND VNB vpwr_clk_buf1_159 vpwr_clk_buf1_159 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_159 VGND VNB vpwr_clk_buf1_159 vpwr_clk_buf1_159 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_160 VGND VNB vpwr_clk_buf1_160 vpwr_clk_buf1_160 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_160 VGND VNB vpwr_clk_buf1_160 vpwr_clk_buf1_160 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_160 VGND VNB vpwr_clk_buf1_160 vpwr_clk_buf1_160 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_161 VGND VNB vpwr_clk_buf1_161 vpwr_clk_buf1_161 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_161 VGND VNB vpwr_clk_buf1_161 vpwr_clk_buf1_161 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_161 VGND VNB vpwr_clk_buf1_161 vpwr_clk_buf1_161 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_162 VGND VNB vpwr_clk_buf1_162 vpwr_clk_buf1_162 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_162 VGND VNB vpwr_clk_buf1_162 vpwr_clk_buf1_162 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_162 VGND VNB vpwr_clk_buf1_162 vpwr_clk_buf1_162 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_163 VGND VNB vpwr_clk_buf1_163 vpwr_clk_buf1_163 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_163 VGND VNB vpwr_clk_buf1_163 vpwr_clk_buf1_163 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_163 VGND VNB vpwr_clk_buf1_163 vpwr_clk_buf1_163 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_164 VGND VNB vpwr_clk_buf1_164 vpwr_clk_buf1_164 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_164 VGND VNB vpwr_clk_buf1_164 vpwr_clk_buf1_164 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_164 VGND VNB vpwr_clk_buf1_164 vpwr_clk_buf1_164 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_165 VGND VNB vpwr_clk_buf1_165 vpwr_clk_buf1_165 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_165 VGND VNB vpwr_clk_buf1_165 vpwr_clk_buf1_165 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_165 VGND VNB vpwr_clk_buf1_165 vpwr_clk_buf1_165 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_166 VGND VNB vpwr_clk_buf1_166 vpwr_clk_buf1_166 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_166 VGND VNB vpwr_clk_buf1_166 vpwr_clk_buf1_166 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_166 VGND VNB vpwr_clk_buf1_166 vpwr_clk_buf1_166 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_167 VGND VNB vpwr_clk_buf1_167 vpwr_clk_buf1_167 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_167 VGND VNB vpwr_clk_buf1_167 vpwr_clk_buf1_167 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_167 VGND VNB vpwr_clk_buf1_167 vpwr_clk_buf1_167 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_168 VGND VNB vpwr_clk_buf1_168 vpwr_clk_buf1_168 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_168 VGND VNB vpwr_clk_buf1_168 vpwr_clk_buf1_168 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_168 VGND VNB vpwr_clk_buf1_168 vpwr_clk_buf1_168 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_169 VGND VNB vpwr_clk_buf1_169 vpwr_clk_buf1_169 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_169 VGND VNB vpwr_clk_buf1_169 vpwr_clk_buf1_169 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_169 VGND VNB vpwr_clk_buf1_169 vpwr_clk_buf1_169 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_170 VGND VNB vpwr_clk_buf1_170 vpwr_clk_buf1_170 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_170 VGND VNB vpwr_clk_buf1_170 vpwr_clk_buf1_170 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_170 VGND VNB vpwr_clk_buf1_170 vpwr_clk_buf1_170 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_171 VGND VNB vpwr_clk_buf1_171 vpwr_clk_buf1_171 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_171 VGND VNB vpwr_clk_buf1_171 vpwr_clk_buf1_171 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_171 VGND VNB vpwr_clk_buf1_171 vpwr_clk_buf1_171 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_172 VGND VNB vpwr_clk_buf1_172 vpwr_clk_buf1_172 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_172 VGND VNB vpwr_clk_buf1_172 vpwr_clk_buf1_172 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_172 VGND VNB vpwr_clk_buf1_172 vpwr_clk_buf1_172 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_173 VGND VNB vpwr_clk_buf1_173 vpwr_clk_buf1_173 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_173 VGND VNB vpwr_clk_buf1_173 vpwr_clk_buf1_173 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_173 VGND VNB vpwr_clk_buf1_173 vpwr_clk_buf1_173 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_174 VGND VNB vpwr_clk_buf1_174 vpwr_clk_buf1_174 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_174 VGND VNB vpwr_clk_buf1_174 vpwr_clk_buf1_174 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_174 VGND VNB vpwr_clk_buf1_174 vpwr_clk_buf1_174 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_175 VGND VNB vpwr_clk_buf1_175 vpwr_clk_buf1_175 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_175 VGND VNB vpwr_clk_buf1_175 vpwr_clk_buf1_175 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_175 VGND VNB vpwr_clk_buf1_175 vpwr_clk_buf1_175 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_176 VGND VNB vpwr_clk_buf1_176 vpwr_clk_buf1_176 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_176 VGND VNB vpwr_clk_buf1_176 vpwr_clk_buf1_176 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_176 VGND VNB vpwr_clk_buf1_176 vpwr_clk_buf1_176 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_177 VGND VNB vpwr_clk_buf1_177 vpwr_clk_buf1_177 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_177 VGND VNB vpwr_clk_buf1_177 vpwr_clk_buf1_177 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_177 VGND VNB vpwr_clk_buf1_177 vpwr_clk_buf1_177 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_178 VGND VNB vpwr_clk_buf1_178 vpwr_clk_buf1_178 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_178 VGND VNB vpwr_clk_buf1_178 vpwr_clk_buf1_178 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_178 VGND VNB vpwr_clk_buf1_178 vpwr_clk_buf1_178 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_179 VGND VNB vpwr_clk_buf1_179 vpwr_clk_buf1_179 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_179 VGND VNB vpwr_clk_buf1_179 vpwr_clk_buf1_179 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_179 VGND VNB vpwr_clk_buf1_179 vpwr_clk_buf1_179 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_180 VGND VNB vpwr_clk_buf1_180 vpwr_clk_buf1_180 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_180 VGND VNB vpwr_clk_buf1_180 vpwr_clk_buf1_180 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_180 VGND VNB vpwr_clk_buf1_180 vpwr_clk_buf1_180 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_181 VGND VNB vpwr_clk_buf1_181 vpwr_clk_buf1_181 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_181 VGND VNB vpwr_clk_buf1_181 vpwr_clk_buf1_181 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_181 VGND VNB vpwr_clk_buf1_181 vpwr_clk_buf1_181 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_182 VGND VNB vpwr_clk_buf1_182 vpwr_clk_buf1_182 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_182 VGND VNB vpwr_clk_buf1_182 vpwr_clk_buf1_182 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_182 VGND VNB vpwr_clk_buf1_182 vpwr_clk_buf1_182 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_183 VGND VNB vpwr_clk_buf1_183 vpwr_clk_buf1_183 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_183 VGND VNB vpwr_clk_buf1_183 vpwr_clk_buf1_183 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_183 VGND VNB vpwr_clk_buf1_183 vpwr_clk_buf1_183 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_184 VGND VNB vpwr_clk_buf1_184 vpwr_clk_buf1_184 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_184 VGND VNB vpwr_clk_buf1_184 vpwr_clk_buf1_184 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_184 VGND VNB vpwr_clk_buf1_184 vpwr_clk_buf1_184 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_185 VGND VNB vpwr_clk_buf1_185 vpwr_clk_buf1_185 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_185 VGND VNB vpwr_clk_buf1_185 vpwr_clk_buf1_185 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_185 VGND VNB vpwr_clk_buf1_185 vpwr_clk_buf1_185 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_186 VGND VNB vpwr_clk_buf1_186 vpwr_clk_buf1_186 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_186 VGND VNB vpwr_clk_buf1_186 vpwr_clk_buf1_186 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_186 VGND VNB vpwr_clk_buf1_186 vpwr_clk_buf1_186 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_187 VGND VNB vpwr_clk_buf1_187 vpwr_clk_buf1_187 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_187 VGND VNB vpwr_clk_buf1_187 vpwr_clk_buf1_187 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_187 VGND VNB vpwr_clk_buf1_187 vpwr_clk_buf1_187 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_188 VGND VNB vpwr_clk_buf1_188 vpwr_clk_buf1_188 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_188 VGND VNB vpwr_clk_buf1_188 vpwr_clk_buf1_188 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_188 VGND VNB vpwr_clk_buf1_188 vpwr_clk_buf1_188 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_189 VGND VNB vpwr_clk_buf1_189 vpwr_clk_buf1_189 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_189 VGND VNB vpwr_clk_buf1_189 vpwr_clk_buf1_189 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_189 VGND VNB vpwr_clk_buf1_189 vpwr_clk_buf1_189 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_190 VGND VNB vpwr_clk_buf1_190 vpwr_clk_buf1_190 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_190 VGND VNB vpwr_clk_buf1_190 vpwr_clk_buf1_190 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_190 VGND VNB vpwr_clk_buf1_190 vpwr_clk_buf1_190 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_191 VGND VNB vpwr_clk_buf1_191 vpwr_clk_buf1_191 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_191 VGND VNB vpwr_clk_buf1_191 vpwr_clk_buf1_191 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_191 VGND VNB vpwr_clk_buf1_191 vpwr_clk_buf1_191 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_192 VGND VNB vpwr_clk_buf1_192 vpwr_clk_buf1_192 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_192 VGND VNB vpwr_clk_buf1_192 vpwr_clk_buf1_192 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_192 VGND VNB vpwr_clk_buf1_192 vpwr_clk_buf1_192 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_193 VGND VNB vpwr_clk_buf1_193 vpwr_clk_buf1_193 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_193 VGND VNB vpwr_clk_buf1_193 vpwr_clk_buf1_193 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_193 VGND VNB vpwr_clk_buf1_193 vpwr_clk_buf1_193 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_194 VGND VNB vpwr_clk_buf1_194 vpwr_clk_buf1_194 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_194 VGND VNB vpwr_clk_buf1_194 vpwr_clk_buf1_194 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_194 VGND VNB vpwr_clk_buf1_194 vpwr_clk_buf1_194 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_195 VGND VNB vpwr_clk_buf1_195 vpwr_clk_buf1_195 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_195 VGND VNB vpwr_clk_buf1_195 vpwr_clk_buf1_195 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_195 VGND VNB vpwr_clk_buf1_195 vpwr_clk_buf1_195 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_196 VGND VNB vpwr_clk_buf1_196 vpwr_clk_buf1_196 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_196 VGND VNB vpwr_clk_buf1_196 vpwr_clk_buf1_196 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_196 VGND VNB vpwr_clk_buf1_196 vpwr_clk_buf1_196 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_197 VGND VNB vpwr_clk_buf1_197 vpwr_clk_buf1_197 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_197 VGND VNB vpwr_clk_buf1_197 vpwr_clk_buf1_197 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_197 VGND VNB vpwr_clk_buf1_197 vpwr_clk_buf1_197 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_198 VGND VNB vpwr_clk_buf1_198 vpwr_clk_buf1_198 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_198 VGND VNB vpwr_clk_buf1_198 vpwr_clk_buf1_198 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_198 VGND VNB vpwr_clk_buf1_198 vpwr_clk_buf1_198 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_199 VGND VNB vpwr_clk_buf1_199 vpwr_clk_buf1_199 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_199 VGND VNB vpwr_clk_buf1_199 vpwr_clk_buf1_199 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_199 VGND VNB vpwr_clk_buf1_199 vpwr_clk_buf1_199 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_200 VGND VNB vpwr_clk_buf1_200 vpwr_clk_buf1_200 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_200 VGND VNB vpwr_clk_buf1_200 vpwr_clk_buf1_200 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_200 VGND VNB vpwr_clk_buf1_200 vpwr_clk_buf1_200 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_201 VGND VNB vpwr_clk_buf1_201 vpwr_clk_buf1_201 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_201 VGND VNB vpwr_clk_buf1_201 vpwr_clk_buf1_201 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_201 VGND VNB vpwr_clk_buf1_201 vpwr_clk_buf1_201 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_202 VGND VNB vpwr_clk_buf1_202 vpwr_clk_buf1_202 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_202 VGND VNB vpwr_clk_buf1_202 vpwr_clk_buf1_202 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_202 VGND VNB vpwr_clk_buf1_202 vpwr_clk_buf1_202 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_203 VGND VNB vpwr_clk_buf1_203 vpwr_clk_buf1_203 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_203 VGND VNB vpwr_clk_buf1_203 vpwr_clk_buf1_203 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_203 VGND VNB vpwr_clk_buf1_203 vpwr_clk_buf1_203 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_204 VGND VNB vpwr_clk_buf1_204 vpwr_clk_buf1_204 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_204 VGND VNB vpwr_clk_buf1_204 vpwr_clk_buf1_204 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_204 VGND VNB vpwr_clk_buf1_204 vpwr_clk_buf1_204 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_205 VGND VNB vpwr_clk_buf1_205 vpwr_clk_buf1_205 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_205 VGND VNB vpwr_clk_buf1_205 vpwr_clk_buf1_205 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_205 VGND VNB vpwr_clk_buf1_205 vpwr_clk_buf1_205 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_206 VGND VNB vpwr_clk_buf1_206 vpwr_clk_buf1_206 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_206 VGND VNB vpwr_clk_buf1_206 vpwr_clk_buf1_206 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_206 VGND VNB vpwr_clk_buf1_206 vpwr_clk_buf1_206 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_207 VGND VNB vpwr_clk_buf1_207 vpwr_clk_buf1_207 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_207 VGND VNB vpwr_clk_buf1_207 vpwr_clk_buf1_207 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_207 VGND VNB vpwr_clk_buf1_207 vpwr_clk_buf1_207 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_208 VGND VNB vpwr_clk_buf1_208 vpwr_clk_buf1_208 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_208 VGND VNB vpwr_clk_buf1_208 vpwr_clk_buf1_208 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_208 VGND VNB vpwr_clk_buf1_208 vpwr_clk_buf1_208 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_209 VGND VNB vpwr_clk_buf1_209 vpwr_clk_buf1_209 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_209 VGND VNB vpwr_clk_buf1_209 vpwr_clk_buf1_209 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_209 VGND VNB vpwr_clk_buf1_209 vpwr_clk_buf1_209 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_210 VGND VNB vpwr_clk_buf1_210 vpwr_clk_buf1_210 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_210 VGND VNB vpwr_clk_buf1_210 vpwr_clk_buf1_210 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_210 VGND VNB vpwr_clk_buf1_210 vpwr_clk_buf1_210 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_211 VGND VNB vpwr_clk_buf1_211 vpwr_clk_buf1_211 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_211 VGND VNB vpwr_clk_buf1_211 vpwr_clk_buf1_211 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_211 VGND VNB vpwr_clk_buf1_211 vpwr_clk_buf1_211 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_212 VGND VNB vpwr_clk_buf1_212 vpwr_clk_buf1_212 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_212 VGND VNB vpwr_clk_buf1_212 vpwr_clk_buf1_212 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_212 VGND VNB vpwr_clk_buf1_212 vpwr_clk_buf1_212 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_213 VGND VNB vpwr_clk_buf1_213 vpwr_clk_buf1_213 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_213 VGND VNB vpwr_clk_buf1_213 vpwr_clk_buf1_213 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_213 VGND VNB vpwr_clk_buf1_213 vpwr_clk_buf1_213 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_214 VGND VNB vpwr_clk_buf1_214 vpwr_clk_buf1_214 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_214 VGND VNB vpwr_clk_buf1_214 vpwr_clk_buf1_214 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_214 VGND VNB vpwr_clk_buf1_214 vpwr_clk_buf1_214 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_215 VGND VNB vpwr_clk_buf1_215 vpwr_clk_buf1_215 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_215 VGND VNB vpwr_clk_buf1_215 vpwr_clk_buf1_215 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_215 VGND VNB vpwr_clk_buf1_215 vpwr_clk_buf1_215 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_216 VGND VNB vpwr_clk_buf1_216 vpwr_clk_buf1_216 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_216 VGND VNB vpwr_clk_buf1_216 vpwr_clk_buf1_216 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_216 VGND VNB vpwr_clk_buf1_216 vpwr_clk_buf1_216 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_217 VGND VNB vpwr_clk_buf1_217 vpwr_clk_buf1_217 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_217 VGND VNB vpwr_clk_buf1_217 vpwr_clk_buf1_217 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_217 VGND VNB vpwr_clk_buf1_217 vpwr_clk_buf1_217 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_218 VGND VNB vpwr_clk_buf1_218 vpwr_clk_buf1_218 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_218 VGND VNB vpwr_clk_buf1_218 vpwr_clk_buf1_218 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_218 VGND VNB vpwr_clk_buf1_218 vpwr_clk_buf1_218 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_219 VGND VNB vpwr_clk_buf1_219 vpwr_clk_buf1_219 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_219 VGND VNB vpwr_clk_buf1_219 vpwr_clk_buf1_219 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_219 VGND VNB vpwr_clk_buf1_219 vpwr_clk_buf1_219 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_220 VGND VNB vpwr_clk_buf1_220 vpwr_clk_buf1_220 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_220 VGND VNB vpwr_clk_buf1_220 vpwr_clk_buf1_220 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_220 VGND VNB vpwr_clk_buf1_220 vpwr_clk_buf1_220 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_221 VGND VNB vpwr_clk_buf1_221 vpwr_clk_buf1_221 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_221 VGND VNB vpwr_clk_buf1_221 vpwr_clk_buf1_221 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_221 VGND VNB vpwr_clk_buf1_221 vpwr_clk_buf1_221 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_222 VGND VNB vpwr_clk_buf1_222 vpwr_clk_buf1_222 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_222 VGND VNB vpwr_clk_buf1_222 vpwr_clk_buf1_222 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_222 VGND VNB vpwr_clk_buf1_222 vpwr_clk_buf1_222 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_223 VGND VNB vpwr_clk_buf1_223 vpwr_clk_buf1_223 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_223 VGND VNB vpwr_clk_buf1_223 vpwr_clk_buf1_223 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_223 VGND VNB vpwr_clk_buf1_223 vpwr_clk_buf1_223 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_224 VGND VNB vpwr_clk_buf1_224 vpwr_clk_buf1_224 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_224 VGND VNB vpwr_clk_buf1_224 vpwr_clk_buf1_224 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_224 VGND VNB vpwr_clk_buf1_224 vpwr_clk_buf1_224 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_225 VGND VNB vpwr_clk_buf1_225 vpwr_clk_buf1_225 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_225 VGND VNB vpwr_clk_buf1_225 vpwr_clk_buf1_225 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_225 VGND VNB vpwr_clk_buf1_225 vpwr_clk_buf1_225 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_226 VGND VNB vpwr_clk_buf1_226 vpwr_clk_buf1_226 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_226 VGND VNB vpwr_clk_buf1_226 vpwr_clk_buf1_226 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_226 VGND VNB vpwr_clk_buf1_226 vpwr_clk_buf1_226 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_227 VGND VNB vpwr_clk_buf1_227 vpwr_clk_buf1_227 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_227 VGND VNB vpwr_clk_buf1_227 vpwr_clk_buf1_227 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_227 VGND VNB vpwr_clk_buf1_227 vpwr_clk_buf1_227 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_228 VGND VNB vpwr_clk_buf1_228 vpwr_clk_buf1_228 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_228 VGND VNB vpwr_clk_buf1_228 vpwr_clk_buf1_228 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_228 VGND VNB vpwr_clk_buf1_228 vpwr_clk_buf1_228 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_229 VGND VNB vpwr_clk_buf1_229 vpwr_clk_buf1_229 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_229 VGND VNB vpwr_clk_buf1_229 vpwr_clk_buf1_229 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_229 VGND VNB vpwr_clk_buf1_229 vpwr_clk_buf1_229 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_230 VGND VNB vpwr_clk_buf1_230 vpwr_clk_buf1_230 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_230 VGND VNB vpwr_clk_buf1_230 vpwr_clk_buf1_230 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_230 VGND VNB vpwr_clk_buf1_230 vpwr_clk_buf1_230 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_231 VGND VNB vpwr_clk_buf1_231 vpwr_clk_buf1_231 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_231 VGND VNB vpwr_clk_buf1_231 vpwr_clk_buf1_231 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_231 VGND VNB vpwr_clk_buf1_231 vpwr_clk_buf1_231 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_232 VGND VNB vpwr_clk_buf1_232 vpwr_clk_buf1_232 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_232 VGND VNB vpwr_clk_buf1_232 vpwr_clk_buf1_232 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_232 VGND VNB vpwr_clk_buf1_232 vpwr_clk_buf1_232 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_233 VGND VNB vpwr_clk_buf1_233 vpwr_clk_buf1_233 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_233 VGND VNB vpwr_clk_buf1_233 vpwr_clk_buf1_233 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_233 VGND VNB vpwr_clk_buf1_233 vpwr_clk_buf1_233 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_234 VGND VNB vpwr_clk_buf1_234 vpwr_clk_buf1_234 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_234 VGND VNB vpwr_clk_buf1_234 vpwr_clk_buf1_234 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_234 VGND VNB vpwr_clk_buf1_234 vpwr_clk_buf1_234 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_235 VGND VNB vpwr_clk_buf1_235 vpwr_clk_buf1_235 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_235 VGND VNB vpwr_clk_buf1_235 vpwr_clk_buf1_235 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_235 VGND VNB vpwr_clk_buf1_235 vpwr_clk_buf1_235 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_236 VGND VNB vpwr_clk_buf1_236 vpwr_clk_buf1_236 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_236 VGND VNB vpwr_clk_buf1_236 vpwr_clk_buf1_236 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_236 VGND VNB vpwr_clk_buf1_236 vpwr_clk_buf1_236 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_237 VGND VNB vpwr_clk_buf1_237 vpwr_clk_buf1_237 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_237 VGND VNB vpwr_clk_buf1_237 vpwr_clk_buf1_237 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_237 VGND VNB vpwr_clk_buf1_237 vpwr_clk_buf1_237 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_238 VGND VNB vpwr_clk_buf1_238 vpwr_clk_buf1_238 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_238 VGND VNB vpwr_clk_buf1_238 vpwr_clk_buf1_238 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_238 VGND VNB vpwr_clk_buf1_238 vpwr_clk_buf1_238 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_239 VGND VNB vpwr_clk_buf1_239 vpwr_clk_buf1_239 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_239 VGND VNB vpwr_clk_buf1_239 vpwr_clk_buf1_239 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_239 VGND VNB vpwr_clk_buf1_239 vpwr_clk_buf1_239 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_240 VGND VNB vpwr_clk_buf1_240 vpwr_clk_buf1_240 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_240 VGND VNB vpwr_clk_buf1_240 vpwr_clk_buf1_240 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_240 VGND VNB vpwr_clk_buf1_240 vpwr_clk_buf1_240 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_241 VGND VNB vpwr_clk_buf1_241 vpwr_clk_buf1_241 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_241 VGND VNB vpwr_clk_buf1_241 vpwr_clk_buf1_241 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_241 VGND VNB vpwr_clk_buf1_241 vpwr_clk_buf1_241 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_242 VGND VNB vpwr_clk_buf1_242 vpwr_clk_buf1_242 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_242 VGND VNB vpwr_clk_buf1_242 vpwr_clk_buf1_242 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_242 VGND VNB vpwr_clk_buf1_242 vpwr_clk_buf1_242 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_243 VGND VNB vpwr_clk_buf1_243 vpwr_clk_buf1_243 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_243 VGND VNB vpwr_clk_buf1_243 vpwr_clk_buf1_243 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_243 VGND VNB vpwr_clk_buf1_243 vpwr_clk_buf1_243 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_244 VGND VNB vpwr_clk_buf1_244 vpwr_clk_buf1_244 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_244 VGND VNB vpwr_clk_buf1_244 vpwr_clk_buf1_244 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_244 VGND VNB vpwr_clk_buf1_244 vpwr_clk_buf1_244 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_245 VGND VNB vpwr_clk_buf1_245 vpwr_clk_buf1_245 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_245 VGND VNB vpwr_clk_buf1_245 vpwr_clk_buf1_245 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_245 VGND VNB vpwr_clk_buf1_245 vpwr_clk_buf1_245 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_246 VGND VNB vpwr_clk_buf1_246 vpwr_clk_buf1_246 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_246 VGND VNB vpwr_clk_buf1_246 vpwr_clk_buf1_246 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_246 VGND VNB vpwr_clk_buf1_246 vpwr_clk_buf1_246 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_247 VGND VNB vpwr_clk_buf1_247 vpwr_clk_buf1_247 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_247 VGND VNB vpwr_clk_buf1_247 vpwr_clk_buf1_247 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_247 VGND VNB vpwr_clk_buf1_247 vpwr_clk_buf1_247 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_248 VGND VNB vpwr_clk_buf1_248 vpwr_clk_buf1_248 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_248 VGND VNB vpwr_clk_buf1_248 vpwr_clk_buf1_248 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_248 VGND VNB vpwr_clk_buf1_248 vpwr_clk_buf1_248 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_249 VGND VNB vpwr_clk_buf1_249 vpwr_clk_buf1_249 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_249 VGND VNB vpwr_clk_buf1_249 vpwr_clk_buf1_249 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_249 VGND VNB vpwr_clk_buf1_249 vpwr_clk_buf1_249 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_250 VGND VNB vpwr_clk_buf1_250 vpwr_clk_buf1_250 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_250 VGND VNB vpwr_clk_buf1_250 vpwr_clk_buf1_250 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_250 VGND VNB vpwr_clk_buf1_250 vpwr_clk_buf1_250 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_251 VGND VNB vpwr_clk_buf1_251 vpwr_clk_buf1_251 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_251 VGND VNB vpwr_clk_buf1_251 vpwr_clk_buf1_251 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_251 VGND VNB vpwr_clk_buf1_251 vpwr_clk_buf1_251 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_252 VGND VNB vpwr_clk_buf1_252 vpwr_clk_buf1_252 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_252 VGND VNB vpwr_clk_buf1_252 vpwr_clk_buf1_252 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_252 VGND VNB vpwr_clk_buf1_252 vpwr_clk_buf1_252 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_253 VGND VNB vpwr_clk_buf1_253 vpwr_clk_buf1_253 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_253 VGND VNB vpwr_clk_buf1_253 vpwr_clk_buf1_253 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_253 VGND VNB vpwr_clk_buf1_253 vpwr_clk_buf1_253 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_254 VGND VNB vpwr_clk_buf1_254 vpwr_clk_buf1_254 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_254 VGND VNB vpwr_clk_buf1_254 vpwr_clk_buf1_254 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_254 VGND VNB vpwr_clk_buf1_254 vpwr_clk_buf1_254 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_255 VGND VNB vpwr_clk_buf1_255 vpwr_clk_buf1_255 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_255 VGND VNB vpwr_clk_buf1_255 vpwr_clk_buf1_255 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_255 VGND VNB vpwr_clk_buf1_255 vpwr_clk_buf1_255 sky130_fd_sc_hd__decap_12

VC_0  clk_0  VGND pulse 0 1.8 1.14n 1n 1n 48n 100n
VC_1  clk_1  VGND pulse 0 1.8  1.0n 1n 1n 48n 100n
VC_2  clk_2  VGND pulse 0 1.8 0.96n 1n 1n 48n 100n
VC_3  clk_3  VGND pulse 0 1.8 0.45n 1n 1n 48n 100n
VC_4  clk_4  VGND pulse 0 1.8 0.81n 1n 1n 48n 100n
VC_5  clk_5  VGND pulse 0 1.8 1.96n 1n 1n 48n 100n
VC_6  clk_6  VGND pulse 0 1.8 1.12n 1n 1n 48n 100n
VC_7  clk_7  VGND pulse 0 1.8 1.11n 1n 1n 48n 100n
VC_8  clk_8  VGND pulse 0 1.8  1.5n 1n 1n 48n 100n
VC_9  clk_9  VGND pulse 0 1.8 0.86n 1n 1n 48n 100n
VC_10 clk_10 VGND pulse 0 1.8  0.6n 1n 1n 48n 100n
VC_11 clk_11 VGND pulse 0 1.8 1.37n 1n 1n 48n 100n
VC_12 clk_12 VGND pulse 0 1.8 1.93n 1n 1n 48n 100n
VC_13 clk_13 VGND pulse 0 1.8 0.84n 1n 1n 48n 100n
VC_14 clk_14 VGND pulse 0 1.8 0.94n 1n 1n 48n 100n
VC_15 clk_15 VGND pulse 0 1.8 0.08n 1n 1n 48n 100n
VC_16 clk_16 VGND pulse 0 1.8 0.54n 1n 1n 48n 100n
VC_17 clk_17 VGND pulse 0 1.8 1.44n 1n 1n 48n 100n
VC_18 clk_18 VGND pulse 0 1.8 0.66n 1n 1n 48n 100n
VC_19 clk_19 VGND pulse 0 1.8 1.05n 1n 1n 48n 100n
VC_20 clk_20 VGND pulse 0 1.8 0.64n 1n 1n 48n 100n
VC_21 clk_21 VGND pulse 0 1.8 1.54n 1n 1n 48n 100n
VC_22 clk_22 VGND pulse 0 1.8 0.19n 1n 1n 48n 100n
VC_23 clk_23 VGND pulse 0 1.8 1.57n 1n 1n 48n 100n
VC_24 clk_24 VGND pulse 0 1.8 1.81n 1n 1n 48n 100n
VC_25 clk_25 VGND pulse 0 1.8 0.61n 1n 1n 48n 100n
VC_26 clk_26 VGND pulse 0 1.8 1.27n 1n 1n 48n 100n
VC_27 clk_27 VGND pulse 0 1.8  1.4n 1n 1n 48n 100n
VC_28 clk_28 VGND pulse 0 1.8 0.86n 1n 1n 48n 100n
VC_29 clk_29 VGND pulse 0 1.8  1.5n 1n 1n 48n 100n
VC_30 clk_30 VGND pulse 0 1.8 1.41n 1n 1n 48n 100n
VC_31 clk_31 VGND pulse 0 1.8 1.05n 1n 1n 48n 100n

x0_0  clk_0  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  co_0  sky130_fd_sc_hd__clkbuf_1
x0_1  clk_1  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  co_1  sky130_fd_sc_hd__clkbuf_1
x0_2  clk_2  VGND VNB vpwr_clk_buf1_2  vpwr_clk_buf1_2  co_2  sky130_fd_sc_hd__clkbuf_1
x0_3  clk_3  VGND VNB vpwr_clk_buf1_3  vpwr_clk_buf1_3  co_3  sky130_fd_sc_hd__clkbuf_1
x0_4  clk_4  VGND VNB vpwr_clk_buf1_4  vpwr_clk_buf1_4  co_4  sky130_fd_sc_hd__clkbuf_1
x0_5  clk_5  VGND VNB vpwr_clk_buf1_5  vpwr_clk_buf1_5  co_5  sky130_fd_sc_hd__clkbuf_1
x0_6  clk_6  VGND VNB vpwr_clk_buf1_6  vpwr_clk_buf1_6  co_6  sky130_fd_sc_hd__clkbuf_1
x0_7  clk_7  VGND VNB vpwr_clk_buf1_7  vpwr_clk_buf1_7  co_7  sky130_fd_sc_hd__clkbuf_1
x0_8  clk_8  VGND VNB vpwr_clk_buf1_8  vpwr_clk_buf1_8  co_8  sky130_fd_sc_hd__clkbuf_1
x0_9  clk_9  VGND VNB vpwr_clk_buf1_9  vpwr_clk_buf1_9  co_9  sky130_fd_sc_hd__clkbuf_1
x0_10 clk_10 VGND VNB vpwr_clk_buf1_10 vpwr_clk_buf1_10 co_10 sky130_fd_sc_hd__clkbuf_1
x0_11 clk_11 VGND VNB vpwr_clk_buf1_11 vpwr_clk_buf1_11 co_11 sky130_fd_sc_hd__clkbuf_1
x0_12 clk_12 VGND VNB vpwr_clk_buf1_12 vpwr_clk_buf1_12 co_12 sky130_fd_sc_hd__clkbuf_1
x0_13 clk_13 VGND VNB vpwr_clk_buf1_13 vpwr_clk_buf1_13 co_13 sky130_fd_sc_hd__clkbuf_1
x0_14 clk_14 VGND VNB vpwr_clk_buf1_14 vpwr_clk_buf1_14 co_14 sky130_fd_sc_hd__clkbuf_1
x0_15 clk_15 VGND VNB vpwr_clk_buf1_15 vpwr_clk_buf1_15 co_15 sky130_fd_sc_hd__clkbuf_1
x0_16 clk_16 VGND VNB vpwr_clk_buf1_16 vpwr_clk_buf1_16 co_16 sky130_fd_sc_hd__clkbuf_1
x0_17 clk_17 VGND VNB vpwr_clk_buf1_17 vpwr_clk_buf1_17 co_17 sky130_fd_sc_hd__clkbuf_1
x0_18 clk_18 VGND VNB vpwr_clk_buf1_18 vpwr_clk_buf1_18 co_18 sky130_fd_sc_hd__clkbuf_1
x0_19 clk_19 VGND VNB vpwr_clk_buf1_19 vpwr_clk_buf1_19 co_19 sky130_fd_sc_hd__clkbuf_1
x0_20 clk_20 VGND VNB vpwr_clk_buf1_20 vpwr_clk_buf1_20 co_20 sky130_fd_sc_hd__clkbuf_1
x0_21 clk_21 VGND VNB vpwr_clk_buf1_21 vpwr_clk_buf1_21 co_21 sky130_fd_sc_hd__clkbuf_1
x0_22 clk_22 VGND VNB vpwr_clk_buf1_22 vpwr_clk_buf1_22 co_22 sky130_fd_sc_hd__clkbuf_1
x0_23 clk_23 VGND VNB vpwr_clk_buf1_23 vpwr_clk_buf1_23 co_23 sky130_fd_sc_hd__clkbuf_1
x0_24 clk_24 VGND VNB vpwr_clk_buf1_24 vpwr_clk_buf1_24 co_24 sky130_fd_sc_hd__clkbuf_1
x0_25 clk_25 VGND VNB vpwr_clk_buf1_25 vpwr_clk_buf1_25 co_25 sky130_fd_sc_hd__clkbuf_1
x0_26 clk_26 VGND VNB vpwr_clk_buf1_26 vpwr_clk_buf1_26 co_26 sky130_fd_sc_hd__clkbuf_1
x0_27 clk_27 VGND VNB vpwr_clk_buf1_27 vpwr_clk_buf1_27 co_27 sky130_fd_sc_hd__clkbuf_1
x0_28 clk_28 VGND VNB vpwr_clk_buf1_28 vpwr_clk_buf1_28 co_28 sky130_fd_sc_hd__clkbuf_1
x0_29 clk_29 VGND VNB vpwr_clk_buf1_29 vpwr_clk_buf1_29 co_29 sky130_fd_sc_hd__clkbuf_1
x0_30 clk_30 VGND VNB vpwr_clk_buf1_30 vpwr_clk_buf1_30 co_30 sky130_fd_sc_hd__clkbuf_1
x0_31 clk_31 VGND VNB vpwr_clk_buf1_31 vpwr_clk_buf1_31 co_31 sky130_fd_sc_hd__clkbuf_1

xdiode_0  co_0  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_1  co_1  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_2  co_2  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_3  co_3  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_4  co_4  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_5  co_5  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_6  co_6  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_7  co_7  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_8  co_8  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_9  co_9  VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_10 co_10 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_11 co_11 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_12 co_12 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_13 co_13 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_14 co_14 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_15 co_15 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_16 co_16 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_17 co_17 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_18 co_18 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_19 co_19 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_20 co_20 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_21 co_21 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_22 co_22 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_23 co_23 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_24 co_24 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_25 co_25 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_26 co_26 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_27 co_27 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_28 co_28 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_29 co_29 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_30 co_30 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2
xdiode_31 co_31 VGND VNB vpwr_0 vpwr_0 sky130_fd_sc_hd__diode_2

R_0  co_0  co_1  ${RLOAD}
R_1  co_1  co_2  ${RLOAD}
R_2  co_2  co_3  ${RLOAD}
R_3  co_3  co_4  ${RLOAD}
R_4  co_4  co_5  ${RLOAD}
R_5  co_5  co_6  ${RLOAD}
R_6  co_6  co_7  ${RLOAD}
R_7  co_7  co_8  ${RLOAD}
R_8  co_8  co_9  ${RLOAD}
R_9  co_9  co_10 ${RLOAD}
R_10 co_10 co_11 ${RLOAD}
R_11 co_11 co_12 ${RLOAD}
R_12 co_12 co_13 ${RLOAD}
R_13 co_13 co_14 ${RLOAD}
R_14 co_14 co_15 ${RLOAD}
R_15 co_15 co_16 ${RLOAD}
R_16 co_16 co_17 ${RLOAD}
R_17 co_17 co_18 ${RLOAD}
R_18 co_18 co_19 ${RLOAD}
R_19 co_19 co_20 ${RLOAD}
R_20 co_20 co_21 ${RLOAD}
R_21 co_21 co_22 ${RLOAD}
R_22 co_22 co_23 ${RLOAD}
R_23 co_23 co_24 ${RLOAD}
R_24 co_24 co_25 ${RLOAD}
R_25 co_25 co_26 ${RLOAD}
R_26 co_26 co_27 ${RLOAD}
R_27 co_27 co_28 ${RLOAD}
R_28 co_28 co_29 ${RLOAD}
R_29 co_29 co_30 ${RLOAD}
R_30 co_30 co_31 ${RLOAD}
R_31 co_31 co_32 ${RLOAD}

x1_0_0  co_0  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0  sky130_fd_sc_hd__clkbuf_16
x1_1_0  co_0  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_0  sky130_fd_sc_hd__clkbuf_16
x1_2_0  co_0  VGND VNB vpwr_clk_buf1_2  vpwr_clk_buf1_2  ff_0  sky130_fd_sc_hd__clkbuf_16
x1_3_0  co_0  VGND VNB vpwr_clk_buf1_3  vpwr_clk_buf1_3  ff_0  sky130_fd_sc_hd__clkbuf_16
x1_4_0  co_0  VGND VNB vpwr_clk_buf1_4  vpwr_clk_buf1_4  ff_0  sky130_fd_sc_hd__clkbuf_16
x1_5_0  co_0  VGND VNB vpwr_clk_buf1_5  vpwr_clk_buf1_5  ff_0  sky130_fd_sc_hd__clkbuf_16
x1_6_0  co_0  VGND VNB vpwr_clk_buf1_6  vpwr_clk_buf1_6  ff_0  sky130_fd_sc_hd__clkbuf_16
x1_7_0  co_0  VGND VNB vpwr_clk_buf1_7  vpwr_clk_buf1_7  ff_0  sky130_fd_sc_hd__clkbuf_16
x1_0_1  co_1  VGND VNB vpwr_clk_buf1_8  vpwr_clk_buf1_8  ff_1  sky130_fd_sc_hd__clkbuf_16
x1_1_1  co_1  VGND VNB vpwr_clk_buf1_9  vpwr_clk_buf1_9  ff_1  sky130_fd_sc_hd__clkbuf_16
x1_2_1  co_1  VGND VNB vpwr_clk_buf1_10 vpwr_clk_buf1_10 ff_1  sky130_fd_sc_hd__clkbuf_16
x1_3_1  co_1  VGND VNB vpwr_clk_buf1_11 vpwr_clk_buf1_11 ff_1  sky130_fd_sc_hd__clkbuf_16
x1_4_1  co_1  VGND VNB vpwr_clk_buf1_12 vpwr_clk_buf1_12 ff_1  sky130_fd_sc_hd__clkbuf_16
x1_5_1  co_1  VGND VNB vpwr_clk_buf1_13 vpwr_clk_buf1_13 ff_1  sky130_fd_sc_hd__clkbuf_16
x1_6_1  co_1  VGND VNB vpwr_clk_buf1_14 vpwr_clk_buf1_14 ff_1  sky130_fd_sc_hd__clkbuf_16
x1_7_1  co_1  VGND VNB vpwr_clk_buf1_15 vpwr_clk_buf1_15 ff_1  sky130_fd_sc_hd__clkbuf_16
x1_0_2  co_2  VGND VNB vpwr_clk_buf1_16 vpwr_clk_buf1_16 ff_2  sky130_fd_sc_hd__clkbuf_16
x1_1_2  co_2  VGND VNB vpwr_clk_buf1_17 vpwr_clk_buf1_17 ff_2  sky130_fd_sc_hd__clkbuf_16
x1_2_2  co_2  VGND VNB vpwr_clk_buf1_18 vpwr_clk_buf1_18 ff_2  sky130_fd_sc_hd__clkbuf_16
x1_3_2  co_2  VGND VNB vpwr_clk_buf1_19 vpwr_clk_buf1_19 ff_2  sky130_fd_sc_hd__clkbuf_16
x1_4_2  co_2  VGND VNB vpwr_clk_buf1_20 vpwr_clk_buf1_20 ff_2  sky130_fd_sc_hd__clkbuf_16
x1_5_2  co_2  VGND VNB vpwr_clk_buf1_21 vpwr_clk_buf1_21 ff_2  sky130_fd_sc_hd__clkbuf_16
x1_6_2  co_2  VGND VNB vpwr_clk_buf1_22 vpwr_clk_buf1_22 ff_2  sky130_fd_sc_hd__clkbuf_16
x1_7_2  co_2  VGND VNB vpwr_clk_buf1_23 vpwr_clk_buf1_23 ff_2  sky130_fd_sc_hd__clkbuf_16
x1_0_3  co_3  VGND VNB vpwr_clk_buf1_24 vpwr_clk_buf1_24 ff_3  sky130_fd_sc_hd__clkbuf_16
x1_1_3  co_3  VGND VNB vpwr_clk_buf1_25 vpwr_clk_buf1_25 ff_3  sky130_fd_sc_hd__clkbuf_16
x1_2_3  co_3  VGND VNB vpwr_clk_buf1_26 vpwr_clk_buf1_26 ff_3  sky130_fd_sc_hd__clkbuf_16
x1_3_3  co_3  VGND VNB vpwr_clk_buf1_27 vpwr_clk_buf1_27 ff_3  sky130_fd_sc_hd__clkbuf_16
x1_4_3  co_3  VGND VNB vpwr_clk_buf1_28 vpwr_clk_buf1_28 ff_3  sky130_fd_sc_hd__clkbuf_16
x1_5_3  co_3  VGND VNB vpwr_clk_buf1_29 vpwr_clk_buf1_29 ff_3  sky130_fd_sc_hd__clkbuf_16
x1_6_3  co_3  VGND VNB vpwr_clk_buf1_30 vpwr_clk_buf1_30 ff_3  sky130_fd_sc_hd__clkbuf_16
x1_7_3  co_3  VGND VNB vpwr_clk_buf1_31 vpwr_clk_buf1_31 ff_3  sky130_fd_sc_hd__clkbuf_16
x1_0_4  co_4  VGND VNB vpwr_clk_buf1_32 vpwr_clk_buf1_32 ff_4  sky130_fd_sc_hd__clkbuf_16
x1_1_4  co_4  VGND VNB vpwr_clk_buf1_33 vpwr_clk_buf1_33 ff_4  sky130_fd_sc_hd__clkbuf_16
x1_2_4  co_4  VGND VNB vpwr_clk_buf1_34 vpwr_clk_buf1_34 ff_4  sky130_fd_sc_hd__clkbuf_16
x1_3_4  co_4  VGND VNB vpwr_clk_buf1_35 vpwr_clk_buf1_35 ff_4  sky130_fd_sc_hd__clkbuf_16
x1_4_4  co_4  VGND VNB vpwr_clk_buf1_36 vpwr_clk_buf1_36 ff_4  sky130_fd_sc_hd__clkbuf_16
x1_5_4  co_4  VGND VNB vpwr_clk_buf1_37 vpwr_clk_buf1_37 ff_4  sky130_fd_sc_hd__clkbuf_16
x1_6_4  co_4  VGND VNB vpwr_clk_buf1_38 vpwr_clk_buf1_38 ff_4  sky130_fd_sc_hd__clkbuf_16
x1_7_4  co_4  VGND VNB vpwr_clk_buf1_39 vpwr_clk_buf1_39 ff_4  sky130_fd_sc_hd__clkbuf_16
x1_0_5  co_5  VGND VNB vpwr_clk_buf1_40 vpwr_clk_buf1_40 ff_5  sky130_fd_sc_hd__clkbuf_16
x1_1_5  co_5  VGND VNB vpwr_clk_buf1_41 vpwr_clk_buf1_41 ff_5  sky130_fd_sc_hd__clkbuf_16
x1_2_5  co_5  VGND VNB vpwr_clk_buf1_42 vpwr_clk_buf1_42 ff_5  sky130_fd_sc_hd__clkbuf_16
x1_3_5  co_5  VGND VNB vpwr_clk_buf1_43 vpwr_clk_buf1_43 ff_5  sky130_fd_sc_hd__clkbuf_16
x1_4_5  co_5  VGND VNB vpwr_clk_buf1_44 vpwr_clk_buf1_44 ff_5  sky130_fd_sc_hd__clkbuf_16
x1_5_5  co_5  VGND VNB vpwr_clk_buf1_45 vpwr_clk_buf1_45 ff_5  sky130_fd_sc_hd__clkbuf_16
x1_6_5  co_5  VGND VNB vpwr_clk_buf1_46 vpwr_clk_buf1_46 ff_5  sky130_fd_sc_hd__clkbuf_16
x1_7_5  co_5  VGND VNB vpwr_clk_buf1_47 vpwr_clk_buf1_47 ff_5  sky130_fd_sc_hd__clkbuf_16
x1_0_6  co_6  VGND VNB vpwr_clk_buf1_48 vpwr_clk_buf1_48 ff_6  sky130_fd_sc_hd__clkbuf_16
x1_1_6  co_6  VGND VNB vpwr_clk_buf1_49 vpwr_clk_buf1_49 ff_6  sky130_fd_sc_hd__clkbuf_16
x1_2_6  co_6  VGND VNB vpwr_clk_buf1_50 vpwr_clk_buf1_50 ff_6  sky130_fd_sc_hd__clkbuf_16
x1_3_6  co_6  VGND VNB vpwr_clk_buf1_51 vpwr_clk_buf1_51 ff_6  sky130_fd_sc_hd__clkbuf_16
x1_4_6  co_6  VGND VNB vpwr_clk_buf1_52 vpwr_clk_buf1_52 ff_6  sky130_fd_sc_hd__clkbuf_16
x1_5_6  co_6  VGND VNB vpwr_clk_buf1_53 vpwr_clk_buf1_53 ff_6  sky130_fd_sc_hd__clkbuf_16
x1_6_6  co_6  VGND VNB vpwr_clk_buf1_54 vpwr_clk_buf1_54 ff_6  sky130_fd_sc_hd__clkbuf_16
x1_7_6  co_6  VGND VNB vpwr_clk_buf1_55 vpwr_clk_buf1_55 ff_6  sky130_fd_sc_hd__clkbuf_16
x1_0_7  co_7  VGND VNB vpwr_clk_buf1_56 vpwr_clk_buf1_56 ff_7  sky130_fd_sc_hd__clkbuf_16
x1_1_7  co_7  VGND VNB vpwr_clk_buf1_57 vpwr_clk_buf1_57 ff_7  sky130_fd_sc_hd__clkbuf_16
x1_2_7  co_7  VGND VNB vpwr_clk_buf1_58 vpwr_clk_buf1_58 ff_7  sky130_fd_sc_hd__clkbuf_16
x1_3_7  co_7  VGND VNB vpwr_clk_buf1_59 vpwr_clk_buf1_59 ff_7  sky130_fd_sc_hd__clkbuf_16
x1_4_7  co_7  VGND VNB vpwr_clk_buf1_60 vpwr_clk_buf1_60 ff_7  sky130_fd_sc_hd__clkbuf_16
x1_5_7  co_7  VGND VNB vpwr_clk_buf1_61 vpwr_clk_buf1_61 ff_7  sky130_fd_sc_hd__clkbuf_16
x1_6_7  co_7  VGND VNB vpwr_clk_buf1_62 vpwr_clk_buf1_62 ff_7  sky130_fd_sc_hd__clkbuf_16
x1_7_7  co_7  VGND VNB vpwr_clk_buf1_63 vpwr_clk_buf1_63 ff_7  sky130_fd_sc_hd__clkbuf_16
x1_0_8  co_8  VGND VNB vpwr_clk_buf1_64 vpwr_clk_buf1_64 ff_8  sky130_fd_sc_hd__clkbuf_16
x1_1_8  co_8  VGND VNB vpwr_clk_buf1_65 vpwr_clk_buf1_65 ff_8  sky130_fd_sc_hd__clkbuf_16
x1_2_8  co_8  VGND VNB vpwr_clk_buf1_66 vpwr_clk_buf1_66 ff_8  sky130_fd_sc_hd__clkbuf_16
x1_3_8  co_8  VGND VNB vpwr_clk_buf1_67 vpwr_clk_buf1_67 ff_8  sky130_fd_sc_hd__clkbuf_16
x1_4_8  co_8  VGND VNB vpwr_clk_buf1_68 vpwr_clk_buf1_68 ff_8  sky130_fd_sc_hd__clkbuf_16
x1_5_8  co_8  VGND VNB vpwr_clk_buf1_69 vpwr_clk_buf1_69 ff_8  sky130_fd_sc_hd__clkbuf_16
x1_6_8  co_8  VGND VNB vpwr_clk_buf1_70 vpwr_clk_buf1_70 ff_8  sky130_fd_sc_hd__clkbuf_16
x1_7_8  co_8  VGND VNB vpwr_clk_buf1_71 vpwr_clk_buf1_71 ff_8  sky130_fd_sc_hd__clkbuf_16
x1_0_9  co_9  VGND VNB vpwr_clk_buf1_72 vpwr_clk_buf1_72 ff_9  sky130_fd_sc_hd__clkbuf_16
x1_1_9  co_9  VGND VNB vpwr_clk_buf1_73 vpwr_clk_buf1_73 ff_9  sky130_fd_sc_hd__clkbuf_16
x1_2_9  co_9  VGND VNB vpwr_clk_buf1_74 vpwr_clk_buf1_74 ff_9  sky130_fd_sc_hd__clkbuf_16
x1_3_9  co_9  VGND VNB vpwr_clk_buf1_75 vpwr_clk_buf1_75 ff_9  sky130_fd_sc_hd__clkbuf_16
x1_4_9  co_9  VGND VNB vpwr_clk_buf1_76 vpwr_clk_buf1_76 ff_9  sky130_fd_sc_hd__clkbuf_16
x1_5_9  co_9  VGND VNB vpwr_clk_buf1_77 vpwr_clk_buf1_77 ff_9  sky130_fd_sc_hd__clkbuf_16
x1_6_9  co_9  VGND VNB vpwr_clk_buf1_78 vpwr_clk_buf1_78 ff_9  sky130_fd_sc_hd__clkbuf_16
x1_7_9  co_9  VGND VNB vpwr_clk_buf1_79 vpwr_clk_buf1_79 ff_9  sky130_fd_sc_hd__clkbuf_16
x1_0_10 co_10 VGND VNB vpwr_clk_buf1_80 vpwr_clk_buf1_80 ff_10 sky130_fd_sc_hd__clkbuf_16
x1_1_10 co_10 VGND VNB vpwr_clk_buf1_81 vpwr_clk_buf1_81 ff_10 sky130_fd_sc_hd__clkbuf_16
x1_2_10 co_10 VGND VNB vpwr_clk_buf1_82 vpwr_clk_buf1_82 ff_10 sky130_fd_sc_hd__clkbuf_16
x1_3_10 co_10 VGND VNB vpwr_clk_buf1_83 vpwr_clk_buf1_83 ff_10 sky130_fd_sc_hd__clkbuf_16
x1_4_10 co_10 VGND VNB vpwr_clk_buf1_84 vpwr_clk_buf1_84 ff_10 sky130_fd_sc_hd__clkbuf_16
x1_5_10 co_10 VGND VNB vpwr_clk_buf1_85 vpwr_clk_buf1_85 ff_10 sky130_fd_sc_hd__clkbuf_16
x1_6_10 co_10 VGND VNB vpwr_clk_buf1_86 vpwr_clk_buf1_86 ff_10 sky130_fd_sc_hd__clkbuf_16
x1_7_10 co_10 VGND VNB vpwr_clk_buf1_87 vpwr_clk_buf1_87 ff_10 sky130_fd_sc_hd__clkbuf_16
x1_0_11 co_11 VGND VNB vpwr_clk_buf1_88 vpwr_clk_buf1_88 ff_11 sky130_fd_sc_hd__clkbuf_16
x1_1_11 co_11 VGND VNB vpwr_clk_buf1_89 vpwr_clk_buf1_89 ff_11 sky130_fd_sc_hd__clkbuf_16
x1_2_11 co_11 VGND VNB vpwr_clk_buf1_90 vpwr_clk_buf1_90 ff_11 sky130_fd_sc_hd__clkbuf_16
x1_3_11 co_11 VGND VNB vpwr_clk_buf1_91 vpwr_clk_buf1_91 ff_11 sky130_fd_sc_hd__clkbuf_16
x1_4_11 co_11 VGND VNB vpwr_clk_buf1_92 vpwr_clk_buf1_92 ff_11 sky130_fd_sc_hd__clkbuf_16
x1_5_11 co_11 VGND VNB vpwr_clk_buf1_93 vpwr_clk_buf1_93 ff_11 sky130_fd_sc_hd__clkbuf_16
x1_6_11 co_11 VGND VNB vpwr_clk_buf1_94 vpwr_clk_buf1_94 ff_11 sky130_fd_sc_hd__clkbuf_16
x1_7_11 co_11 VGND VNB vpwr_clk_buf1_95 vpwr_clk_buf1_95 ff_11 sky130_fd_sc_hd__clkbuf_16
x1_0_12 co_12 VGND VNB vpwr_clk_buf1_96 vpwr_clk_buf1_96 ff_12 sky130_fd_sc_hd__clkbuf_16
x1_1_12 co_12 VGND VNB vpwr_clk_buf1_97 vpwr_clk_buf1_97 ff_12 sky130_fd_sc_hd__clkbuf_16
x1_2_12 co_12 VGND VNB vpwr_clk_buf1_98 vpwr_clk_buf1_98 ff_12 sky130_fd_sc_hd__clkbuf_16
x1_3_12 co_12 VGND VNB vpwr_clk_buf1_99 vpwr_clk_buf1_99 ff_12 sky130_fd_sc_hd__clkbuf_16
x1_4_12 co_12 VGND VNB vpwr_clk_buf1_100 vpwr_clk_buf1_100 ff_12 sky130_fd_sc_hd__clkbuf_16
x1_5_12 co_12 VGND VNB vpwr_clk_buf1_101 vpwr_clk_buf1_101 ff_12 sky130_fd_sc_hd__clkbuf_16
x1_6_12 co_12 VGND VNB vpwr_clk_buf1_102 vpwr_clk_buf1_102 ff_12 sky130_fd_sc_hd__clkbuf_16
x1_7_12 co_12 VGND VNB vpwr_clk_buf1_103 vpwr_clk_buf1_103 ff_12 sky130_fd_sc_hd__clkbuf_16
x1_0_13 co_13 VGND VNB vpwr_clk_buf1_104 vpwr_clk_buf1_104 ff_13 sky130_fd_sc_hd__clkbuf_16
x1_1_13 co_13 VGND VNB vpwr_clk_buf1_105 vpwr_clk_buf1_105 ff_13 sky130_fd_sc_hd__clkbuf_16
x1_2_13 co_13 VGND VNB vpwr_clk_buf1_106 vpwr_clk_buf1_106 ff_13 sky130_fd_sc_hd__clkbuf_16
x1_3_13 co_13 VGND VNB vpwr_clk_buf1_107 vpwr_clk_buf1_107 ff_13 sky130_fd_sc_hd__clkbuf_16
x1_4_13 co_13 VGND VNB vpwr_clk_buf1_108 vpwr_clk_buf1_108 ff_13 sky130_fd_sc_hd__clkbuf_16
x1_5_13 co_13 VGND VNB vpwr_clk_buf1_109 vpwr_clk_buf1_109 ff_13 sky130_fd_sc_hd__clkbuf_16
x1_6_13 co_13 VGND VNB vpwr_clk_buf1_110 vpwr_clk_buf1_110 ff_13 sky130_fd_sc_hd__clkbuf_16
x1_7_13 co_13 VGND VNB vpwr_clk_buf1_111 vpwr_clk_buf1_111 ff_13 sky130_fd_sc_hd__clkbuf_16
x1_0_14 co_14 VGND VNB vpwr_clk_buf1_112 vpwr_clk_buf1_112 ff_14 sky130_fd_sc_hd__clkbuf_16
x1_1_14 co_14 VGND VNB vpwr_clk_buf1_113 vpwr_clk_buf1_113 ff_14 sky130_fd_sc_hd__clkbuf_16
x1_2_14 co_14 VGND VNB vpwr_clk_buf1_114 vpwr_clk_buf1_114 ff_14 sky130_fd_sc_hd__clkbuf_16
x1_3_14 co_14 VGND VNB vpwr_clk_buf1_115 vpwr_clk_buf1_115 ff_14 sky130_fd_sc_hd__clkbuf_16
x1_4_14 co_14 VGND VNB vpwr_clk_buf1_116 vpwr_clk_buf1_116 ff_14 sky130_fd_sc_hd__clkbuf_16
x1_5_14 co_14 VGND VNB vpwr_clk_buf1_117 vpwr_clk_buf1_117 ff_14 sky130_fd_sc_hd__clkbuf_16
x1_6_14 co_14 VGND VNB vpwr_clk_buf1_118 vpwr_clk_buf1_118 ff_14 sky130_fd_sc_hd__clkbuf_16
x1_7_14 co_14 VGND VNB vpwr_clk_buf1_119 vpwr_clk_buf1_119 ff_14 sky130_fd_sc_hd__clkbuf_16
x1_0_15 co_15 VGND VNB vpwr_clk_buf1_120 vpwr_clk_buf1_120 ff_15 sky130_fd_sc_hd__clkbuf_16
x1_1_15 co_15 VGND VNB vpwr_clk_buf1_121 vpwr_clk_buf1_121 ff_15 sky130_fd_sc_hd__clkbuf_16
x1_2_15 co_15 VGND VNB vpwr_clk_buf1_122 vpwr_clk_buf1_122 ff_15 sky130_fd_sc_hd__clkbuf_16
x1_3_15 co_15 VGND VNB vpwr_clk_buf1_123 vpwr_clk_buf1_123 ff_15 sky130_fd_sc_hd__clkbuf_16
x1_4_15 co_15 VGND VNB vpwr_clk_buf1_124 vpwr_clk_buf1_124 ff_15 sky130_fd_sc_hd__clkbuf_16
x1_5_15 co_15 VGND VNB vpwr_clk_buf1_125 vpwr_clk_buf1_125 ff_15 sky130_fd_sc_hd__clkbuf_16
x1_6_15 co_15 VGND VNB vpwr_clk_buf1_126 vpwr_clk_buf1_126 ff_15 sky130_fd_sc_hd__clkbuf_16
x1_7_15 co_15 VGND VNB vpwr_clk_buf1_127 vpwr_clk_buf1_127 ff_15 sky130_fd_sc_hd__clkbuf_16
x1_0_16 co_16 VGND VNB vpwr_clk_buf1_128 vpwr_clk_buf1_128 ff_16 sky130_fd_sc_hd__clkbuf_16
x1_1_16 co_16 VGND VNB vpwr_clk_buf1_129 vpwr_clk_buf1_129 ff_16 sky130_fd_sc_hd__clkbuf_16
x1_2_16 co_16 VGND VNB vpwr_clk_buf1_130 vpwr_clk_buf1_130 ff_16 sky130_fd_sc_hd__clkbuf_16
x1_3_16 co_16 VGND VNB vpwr_clk_buf1_131 vpwr_clk_buf1_131 ff_16 sky130_fd_sc_hd__clkbuf_16
x1_4_16 co_16 VGND VNB vpwr_clk_buf1_132 vpwr_clk_buf1_132 ff_16 sky130_fd_sc_hd__clkbuf_16
x1_5_16 co_16 VGND VNB vpwr_clk_buf1_133 vpwr_clk_buf1_133 ff_16 sky130_fd_sc_hd__clkbuf_16
x1_6_16 co_16 VGND VNB vpwr_clk_buf1_134 vpwr_clk_buf1_134 ff_16 sky130_fd_sc_hd__clkbuf_16
x1_7_16 co_16 VGND VNB vpwr_clk_buf1_135 vpwr_clk_buf1_135 ff_16 sky130_fd_sc_hd__clkbuf_16
x1_0_17 co_17 VGND VNB vpwr_clk_buf1_136 vpwr_clk_buf1_136 ff_17 sky130_fd_sc_hd__clkbuf_16
x1_1_17 co_17 VGND VNB vpwr_clk_buf1_137 vpwr_clk_buf1_137 ff_17 sky130_fd_sc_hd__clkbuf_16
x1_2_17 co_17 VGND VNB vpwr_clk_buf1_138 vpwr_clk_buf1_138 ff_17 sky130_fd_sc_hd__clkbuf_16
x1_3_17 co_17 VGND VNB vpwr_clk_buf1_139 vpwr_clk_buf1_139 ff_17 sky130_fd_sc_hd__clkbuf_16
x1_4_17 co_17 VGND VNB vpwr_clk_buf1_140 vpwr_clk_buf1_140 ff_17 sky130_fd_sc_hd__clkbuf_16
x1_5_17 co_17 VGND VNB vpwr_clk_buf1_141 vpwr_clk_buf1_141 ff_17 sky130_fd_sc_hd__clkbuf_16
x1_6_17 co_17 VGND VNB vpwr_clk_buf1_142 vpwr_clk_buf1_142 ff_17 sky130_fd_sc_hd__clkbuf_16
x1_7_17 co_17 VGND VNB vpwr_clk_buf1_143 vpwr_clk_buf1_143 ff_17 sky130_fd_sc_hd__clkbuf_16
x1_0_18 co_18 VGND VNB vpwr_clk_buf1_144 vpwr_clk_buf1_144 ff_18 sky130_fd_sc_hd__clkbuf_16
x1_1_18 co_18 VGND VNB vpwr_clk_buf1_145 vpwr_clk_buf1_145 ff_18 sky130_fd_sc_hd__clkbuf_16
x1_2_18 co_18 VGND VNB vpwr_clk_buf1_146 vpwr_clk_buf1_146 ff_18 sky130_fd_sc_hd__clkbuf_16
x1_3_18 co_18 VGND VNB vpwr_clk_buf1_147 vpwr_clk_buf1_147 ff_18 sky130_fd_sc_hd__clkbuf_16
x1_4_18 co_18 VGND VNB vpwr_clk_buf1_148 vpwr_clk_buf1_148 ff_18 sky130_fd_sc_hd__clkbuf_16
x1_5_18 co_18 VGND VNB vpwr_clk_buf1_149 vpwr_clk_buf1_149 ff_18 sky130_fd_sc_hd__clkbuf_16
x1_6_18 co_18 VGND VNB vpwr_clk_buf1_150 vpwr_clk_buf1_150 ff_18 sky130_fd_sc_hd__clkbuf_16
x1_7_18 co_18 VGND VNB vpwr_clk_buf1_151 vpwr_clk_buf1_151 ff_18 sky130_fd_sc_hd__clkbuf_16
x1_0_19 co_19 VGND VNB vpwr_clk_buf1_152 vpwr_clk_buf1_152 ff_19 sky130_fd_sc_hd__clkbuf_16
x1_1_19 co_19 VGND VNB vpwr_clk_buf1_153 vpwr_clk_buf1_153 ff_19 sky130_fd_sc_hd__clkbuf_16
x1_2_19 co_19 VGND VNB vpwr_clk_buf1_154 vpwr_clk_buf1_154 ff_19 sky130_fd_sc_hd__clkbuf_16
x1_3_19 co_19 VGND VNB vpwr_clk_buf1_155 vpwr_clk_buf1_155 ff_19 sky130_fd_sc_hd__clkbuf_16
x1_4_19 co_19 VGND VNB vpwr_clk_buf1_156 vpwr_clk_buf1_156 ff_19 sky130_fd_sc_hd__clkbuf_16
x1_5_19 co_19 VGND VNB vpwr_clk_buf1_157 vpwr_clk_buf1_157 ff_19 sky130_fd_sc_hd__clkbuf_16
x1_6_19 co_19 VGND VNB vpwr_clk_buf1_158 vpwr_clk_buf1_158 ff_19 sky130_fd_sc_hd__clkbuf_16
x1_7_19 co_19 VGND VNB vpwr_clk_buf1_159 vpwr_clk_buf1_159 ff_19 sky130_fd_sc_hd__clkbuf_16
x1_0_20 co_20 VGND VNB vpwr_clk_buf1_160 vpwr_clk_buf1_160 ff_20 sky130_fd_sc_hd__clkbuf_16
x1_1_20 co_20 VGND VNB vpwr_clk_buf1_161 vpwr_clk_buf1_161 ff_20 sky130_fd_sc_hd__clkbuf_16
x1_2_20 co_20 VGND VNB vpwr_clk_buf1_162 vpwr_clk_buf1_162 ff_20 sky130_fd_sc_hd__clkbuf_16
x1_3_20 co_20 VGND VNB vpwr_clk_buf1_163 vpwr_clk_buf1_163 ff_20 sky130_fd_sc_hd__clkbuf_16
x1_4_20 co_20 VGND VNB vpwr_clk_buf1_164 vpwr_clk_buf1_164 ff_20 sky130_fd_sc_hd__clkbuf_16
x1_5_20 co_20 VGND VNB vpwr_clk_buf1_165 vpwr_clk_buf1_165 ff_20 sky130_fd_sc_hd__clkbuf_16
x1_6_20 co_20 VGND VNB vpwr_clk_buf1_166 vpwr_clk_buf1_166 ff_20 sky130_fd_sc_hd__clkbuf_16
x1_7_20 co_20 VGND VNB vpwr_clk_buf1_167 vpwr_clk_buf1_167 ff_20 sky130_fd_sc_hd__clkbuf_16
x1_0_21 co_21 VGND VNB vpwr_clk_buf1_168 vpwr_clk_buf1_168 ff_21 sky130_fd_sc_hd__clkbuf_16
x1_1_21 co_21 VGND VNB vpwr_clk_buf1_169 vpwr_clk_buf1_169 ff_21 sky130_fd_sc_hd__clkbuf_16
x1_2_21 co_21 VGND VNB vpwr_clk_buf1_170 vpwr_clk_buf1_170 ff_21 sky130_fd_sc_hd__clkbuf_16
x1_3_21 co_21 VGND VNB vpwr_clk_buf1_171 vpwr_clk_buf1_171 ff_21 sky130_fd_sc_hd__clkbuf_16
x1_4_21 co_21 VGND VNB vpwr_clk_buf1_172 vpwr_clk_buf1_172 ff_21 sky130_fd_sc_hd__clkbuf_16
x1_5_21 co_21 VGND VNB vpwr_clk_buf1_173 vpwr_clk_buf1_173 ff_21 sky130_fd_sc_hd__clkbuf_16
x1_6_21 co_21 VGND VNB vpwr_clk_buf1_174 vpwr_clk_buf1_174 ff_21 sky130_fd_sc_hd__clkbuf_16
x1_7_21 co_21 VGND VNB vpwr_clk_buf1_175 vpwr_clk_buf1_175 ff_21 sky130_fd_sc_hd__clkbuf_16
x1_0_22 co_22 VGND VNB vpwr_clk_buf1_176 vpwr_clk_buf1_176 ff_22 sky130_fd_sc_hd__clkbuf_16
x1_1_22 co_22 VGND VNB vpwr_clk_buf1_177 vpwr_clk_buf1_177 ff_22 sky130_fd_sc_hd__clkbuf_16
x1_2_22 co_22 VGND VNB vpwr_clk_buf1_178 vpwr_clk_buf1_178 ff_22 sky130_fd_sc_hd__clkbuf_16
x1_3_22 co_22 VGND VNB vpwr_clk_buf1_179 vpwr_clk_buf1_179 ff_22 sky130_fd_sc_hd__clkbuf_16
x1_4_22 co_22 VGND VNB vpwr_clk_buf1_180 vpwr_clk_buf1_180 ff_22 sky130_fd_sc_hd__clkbuf_16
x1_5_22 co_22 VGND VNB vpwr_clk_buf1_181 vpwr_clk_buf1_181 ff_22 sky130_fd_sc_hd__clkbuf_16
x1_6_22 co_22 VGND VNB vpwr_clk_buf1_182 vpwr_clk_buf1_182 ff_22 sky130_fd_sc_hd__clkbuf_16
x1_7_22 co_22 VGND VNB vpwr_clk_buf1_183 vpwr_clk_buf1_183 ff_22 sky130_fd_sc_hd__clkbuf_16
x1_0_23 co_23 VGND VNB vpwr_clk_buf1_184 vpwr_clk_buf1_184 ff_23 sky130_fd_sc_hd__clkbuf_16
x1_1_23 co_23 VGND VNB vpwr_clk_buf1_185 vpwr_clk_buf1_185 ff_23 sky130_fd_sc_hd__clkbuf_16
x1_2_23 co_23 VGND VNB vpwr_clk_buf1_186 vpwr_clk_buf1_186 ff_23 sky130_fd_sc_hd__clkbuf_16
x1_3_23 co_23 VGND VNB vpwr_clk_buf1_187 vpwr_clk_buf1_187 ff_23 sky130_fd_sc_hd__clkbuf_16
x1_4_23 co_23 VGND VNB vpwr_clk_buf1_188 vpwr_clk_buf1_188 ff_23 sky130_fd_sc_hd__clkbuf_16
x1_5_23 co_23 VGND VNB vpwr_clk_buf1_189 vpwr_clk_buf1_189 ff_23 sky130_fd_sc_hd__clkbuf_16
x1_6_23 co_23 VGND VNB vpwr_clk_buf1_190 vpwr_clk_buf1_190 ff_23 sky130_fd_sc_hd__clkbuf_16
x1_7_23 co_23 VGND VNB vpwr_clk_buf1_191 vpwr_clk_buf1_191 ff_23 sky130_fd_sc_hd__clkbuf_16
x1_0_24 co_24 VGND VNB vpwr_clk_buf1_192 vpwr_clk_buf1_192 ff_24 sky130_fd_sc_hd__clkbuf_16
x1_1_24 co_24 VGND VNB vpwr_clk_buf1_193 vpwr_clk_buf1_193 ff_24 sky130_fd_sc_hd__clkbuf_16
x1_2_24 co_24 VGND VNB vpwr_clk_buf1_194 vpwr_clk_buf1_194 ff_24 sky130_fd_sc_hd__clkbuf_16
x1_3_24 co_24 VGND VNB vpwr_clk_buf1_195 vpwr_clk_buf1_195 ff_24 sky130_fd_sc_hd__clkbuf_16
x1_4_24 co_24 VGND VNB vpwr_clk_buf1_196 vpwr_clk_buf1_196 ff_24 sky130_fd_sc_hd__clkbuf_16
x1_5_24 co_24 VGND VNB vpwr_clk_buf1_197 vpwr_clk_buf1_197 ff_24 sky130_fd_sc_hd__clkbuf_16
x1_6_24 co_24 VGND VNB vpwr_clk_buf1_198 vpwr_clk_buf1_198 ff_24 sky130_fd_sc_hd__clkbuf_16
x1_7_24 co_24 VGND VNB vpwr_clk_buf1_199 vpwr_clk_buf1_199 ff_24 sky130_fd_sc_hd__clkbuf_16
x1_0_25 co_25 VGND VNB vpwr_clk_buf1_200 vpwr_clk_buf1_200 ff_25 sky130_fd_sc_hd__clkbuf_16
x1_1_25 co_25 VGND VNB vpwr_clk_buf1_201 vpwr_clk_buf1_201 ff_25 sky130_fd_sc_hd__clkbuf_16
x1_2_25 co_25 VGND VNB vpwr_clk_buf1_202 vpwr_clk_buf1_202 ff_25 sky130_fd_sc_hd__clkbuf_16
x1_3_25 co_25 VGND VNB vpwr_clk_buf1_203 vpwr_clk_buf1_203 ff_25 sky130_fd_sc_hd__clkbuf_16
x1_4_25 co_25 VGND VNB vpwr_clk_buf1_204 vpwr_clk_buf1_204 ff_25 sky130_fd_sc_hd__clkbuf_16
x1_5_25 co_25 VGND VNB vpwr_clk_buf1_205 vpwr_clk_buf1_205 ff_25 sky130_fd_sc_hd__clkbuf_16
x1_6_25 co_25 VGND VNB vpwr_clk_buf1_206 vpwr_clk_buf1_206 ff_25 sky130_fd_sc_hd__clkbuf_16
x1_7_25 co_25 VGND VNB vpwr_clk_buf1_207 vpwr_clk_buf1_207 ff_25 sky130_fd_sc_hd__clkbuf_16
x1_0_26 co_26 VGND VNB vpwr_clk_buf1_208 vpwr_clk_buf1_208 ff_26 sky130_fd_sc_hd__clkbuf_16
x1_1_26 co_26 VGND VNB vpwr_clk_buf1_209 vpwr_clk_buf1_209 ff_26 sky130_fd_sc_hd__clkbuf_16
x1_2_26 co_26 VGND VNB vpwr_clk_buf1_210 vpwr_clk_buf1_210 ff_26 sky130_fd_sc_hd__clkbuf_16
x1_3_26 co_26 VGND VNB vpwr_clk_buf1_211 vpwr_clk_buf1_211 ff_26 sky130_fd_sc_hd__clkbuf_16
x1_4_26 co_26 VGND VNB vpwr_clk_buf1_212 vpwr_clk_buf1_212 ff_26 sky130_fd_sc_hd__clkbuf_16
x1_5_26 co_26 VGND VNB vpwr_clk_buf1_213 vpwr_clk_buf1_213 ff_26 sky130_fd_sc_hd__clkbuf_16
x1_6_26 co_26 VGND VNB vpwr_clk_buf1_214 vpwr_clk_buf1_214 ff_26 sky130_fd_sc_hd__clkbuf_16
x1_7_26 co_26 VGND VNB vpwr_clk_buf1_215 vpwr_clk_buf1_215 ff_26 sky130_fd_sc_hd__clkbuf_16
x1_0_27 co_27 VGND VNB vpwr_clk_buf1_216 vpwr_clk_buf1_216 ff_27 sky130_fd_sc_hd__clkbuf_16
x1_1_27 co_27 VGND VNB vpwr_clk_buf1_217 vpwr_clk_buf1_217 ff_27 sky130_fd_sc_hd__clkbuf_16
x1_2_27 co_27 VGND VNB vpwr_clk_buf1_218 vpwr_clk_buf1_218 ff_27 sky130_fd_sc_hd__clkbuf_16
x1_3_27 co_27 VGND VNB vpwr_clk_buf1_219 vpwr_clk_buf1_219 ff_27 sky130_fd_sc_hd__clkbuf_16
x1_4_27 co_27 VGND VNB vpwr_clk_buf1_220 vpwr_clk_buf1_220 ff_27 sky130_fd_sc_hd__clkbuf_16
x1_5_27 co_27 VGND VNB vpwr_clk_buf1_221 vpwr_clk_buf1_221 ff_27 sky130_fd_sc_hd__clkbuf_16
x1_6_27 co_27 VGND VNB vpwr_clk_buf1_222 vpwr_clk_buf1_222 ff_27 sky130_fd_sc_hd__clkbuf_16
x1_7_27 co_27 VGND VNB vpwr_clk_buf1_223 vpwr_clk_buf1_223 ff_27 sky130_fd_sc_hd__clkbuf_16
x1_0_28 co_28 VGND VNB vpwr_clk_buf1_224 vpwr_clk_buf1_224 ff_28 sky130_fd_sc_hd__clkbuf_16
x1_1_28 co_28 VGND VNB vpwr_clk_buf1_225 vpwr_clk_buf1_225 ff_28 sky130_fd_sc_hd__clkbuf_16
x1_2_28 co_28 VGND VNB vpwr_clk_buf1_226 vpwr_clk_buf1_226 ff_28 sky130_fd_sc_hd__clkbuf_16
x1_3_28 co_28 VGND VNB vpwr_clk_buf1_227 vpwr_clk_buf1_227 ff_28 sky130_fd_sc_hd__clkbuf_16
x1_4_28 co_28 VGND VNB vpwr_clk_buf1_228 vpwr_clk_buf1_228 ff_28 sky130_fd_sc_hd__clkbuf_16
x1_5_28 co_28 VGND VNB vpwr_clk_buf1_229 vpwr_clk_buf1_229 ff_28 sky130_fd_sc_hd__clkbuf_16
x1_6_28 co_28 VGND VNB vpwr_clk_buf1_230 vpwr_clk_buf1_230 ff_28 sky130_fd_sc_hd__clkbuf_16
x1_7_28 co_28 VGND VNB vpwr_clk_buf1_231 vpwr_clk_buf1_231 ff_28 sky130_fd_sc_hd__clkbuf_16
x1_0_29 co_29 VGND VNB vpwr_clk_buf1_232 vpwr_clk_buf1_232 ff_29 sky130_fd_sc_hd__clkbuf_16
x1_1_29 co_29 VGND VNB vpwr_clk_buf1_233 vpwr_clk_buf1_233 ff_29 sky130_fd_sc_hd__clkbuf_16
x1_2_29 co_29 VGND VNB vpwr_clk_buf1_234 vpwr_clk_buf1_234 ff_29 sky130_fd_sc_hd__clkbuf_16
x1_3_29 co_29 VGND VNB vpwr_clk_buf1_235 vpwr_clk_buf1_235 ff_29 sky130_fd_sc_hd__clkbuf_16
x1_4_29 co_29 VGND VNB vpwr_clk_buf1_236 vpwr_clk_buf1_236 ff_29 sky130_fd_sc_hd__clkbuf_16
x1_5_29 co_29 VGND VNB vpwr_clk_buf1_237 vpwr_clk_buf1_237 ff_29 sky130_fd_sc_hd__clkbuf_16
x1_6_29 co_29 VGND VNB vpwr_clk_buf1_238 vpwr_clk_buf1_238 ff_29 sky130_fd_sc_hd__clkbuf_16
x1_7_29 co_29 VGND VNB vpwr_clk_buf1_239 vpwr_clk_buf1_239 ff_29 sky130_fd_sc_hd__clkbuf_16
x1_0_30 co_30 VGND VNB vpwr_clk_buf1_240 vpwr_clk_buf1_240 ff_30 sky130_fd_sc_hd__clkbuf_16
x1_1_30 co_30 VGND VNB vpwr_clk_buf1_241 vpwr_clk_buf1_241 ff_30 sky130_fd_sc_hd__clkbuf_16
x1_2_30 co_30 VGND VNB vpwr_clk_buf1_242 vpwr_clk_buf1_242 ff_30 sky130_fd_sc_hd__clkbuf_16
x1_3_30 co_30 VGND VNB vpwr_clk_buf1_243 vpwr_clk_buf1_243 ff_30 sky130_fd_sc_hd__clkbuf_16
x1_4_30 co_30 VGND VNB vpwr_clk_buf1_244 vpwr_clk_buf1_244 ff_30 sky130_fd_sc_hd__clkbuf_16
x1_5_30 co_30 VGND VNB vpwr_clk_buf1_245 vpwr_clk_buf1_245 ff_30 sky130_fd_sc_hd__clkbuf_16
x1_6_30 co_30 VGND VNB vpwr_clk_buf1_246 vpwr_clk_buf1_246 ff_30 sky130_fd_sc_hd__clkbuf_16
x1_7_30 co_30 VGND VNB vpwr_clk_buf1_247 vpwr_clk_buf1_247 ff_30 sky130_fd_sc_hd__clkbuf_16
x1_0_31 co_31 VGND VNB vpwr_clk_buf1_248 vpwr_clk_buf1_248 ff_31 sky130_fd_sc_hd__clkbuf_16
x1_1_31 co_31 VGND VNB vpwr_clk_buf1_249 vpwr_clk_buf1_249 ff_31 sky130_fd_sc_hd__clkbuf_16
x1_2_31 co_31 VGND VNB vpwr_clk_buf1_250 vpwr_clk_buf1_250 ff_31 sky130_fd_sc_hd__clkbuf_16
x1_3_31 co_31 VGND VNB vpwr_clk_buf1_251 vpwr_clk_buf1_251 ff_31 sky130_fd_sc_hd__clkbuf_16
x1_4_31 co_31 VGND VNB vpwr_clk_buf1_252 vpwr_clk_buf1_252 ff_31 sky130_fd_sc_hd__clkbuf_16
x1_5_31 co_31 VGND VNB vpwr_clk_buf1_253 vpwr_clk_buf1_253 ff_31 sky130_fd_sc_hd__clkbuf_16
x1_6_31 co_31 VGND VNB vpwr_clk_buf1_254 vpwr_clk_buf1_254 ff_31 sky130_fd_sc_hd__clkbuf_16
x1_7_31 co_31 VGND VNB vpwr_clk_buf1_255 vpwr_clk_buf1_255 ff_31 sky130_fd_sc_hd__clkbuf_16

X10F_0  vpwr_0 VGND ff_0  Q1   Q2   Q3   Q4   Q5   Q6   Q7   Q8   Q9   Q10   DFXTP_2_10X
X10F_1  vpwr_0 VGND ff_1  Q11  Q12  Q13  Q14  Q15  Q16  Q17  Q18  Q19  Q20   DFXTP_2_10X
X10F_2  vpwr_0 VGND ff_2  Q21  Q22  Q23  Q24  Q25  Q26  Q27  Q28  Q29  Q30   DFXTP_2_10X
X10F_3  vpwr_0 VGND ff_3  Q31  Q32  Q33  Q34  Q35  Q36  Q37  Q38  Q39  Q40   DFXTP_2_10X
X10F_4  vpwr_0 VGND ff_4  Q41  Q42  Q43  Q44  Q45  Q46  Q47  Q48  Q49  Q50   DFXTP_2_10X
X10F_5  vpwr_0 VGND ff_5  Q51  Q52  Q53  Q54  Q55  Q56  Q57  Q58  Q59  Q60   DFXTP_2_10X
X10F_6  vpwr_0 VGND ff_6  Q61  Q62  Q63  Q64  Q65  Q66  Q67  Q68  Q69  Q70   DFXTP_2_10X
X10F_7  vpwr_0 VGND ff_7  Q71  Q72  Q73  Q74  Q75  Q76  Q77  Q78  Q79  Q80   DFXTP_2_10X
X10F_8  vpwr_0 VGND ff_8  Q81  Q82  Q83  Q84  Q85  Q86  Q87  Q88  Q89  Q90   DFXTP_2_10X
X10F_9  vpwr_0 VGND ff_9  Q91  Q92  Q93  Q94  Q95  Q96  Q97  Q98  Q99  Q100  DFXTP_2_10X
X10F_10 vpwr_0 VGND ff_10 Q101 Q102 Q103 Q104 Q105 Q106 Q107 Q108 Q109 Q110  DFXTP_2_10X
X10F_11 vpwr_0 VGND ff_11 Q111 Q112 Q113 Q114 Q115 Q116 Q117 Q118 Q119 Q120  DFXTP_2_10X
X10F_12 vpwr_0 VGND ff_12 Q121 Q122 Q123 Q124 Q125 Q126 Q127 Q128 Q129 Q130  DFXTP_2_10X
X10F_13 vpwr_0 VGND ff_13 Q131 Q132 Q133 Q134 Q135 Q136 Q137 Q138 Q139 Q140  DFXTP_2_10X
X10F_14 vpwr_0 VGND ff_14 Q141 Q142 Q143 Q144 Q145 Q146 Q147 Q148 Q149 Q150  DFXTP_2_10X
X10F_15 vpwr_0 VGND ff_15 Q151 Q152 Q153 Q154 Q155 Q156 Q157 Q158 Q159 Q160  DFXTP_2_10X
X10F_16 vpwr_0 VGND ff_16 Q161 Q162 Q163 Q164 Q165 Q166 Q167 Q168 Q169 Q170  DFXTP_2_10X
X10F_17 vpwr_0 VGND ff_17 Q171 Q172 Q173 Q174 Q175 Q176 Q177 Q178 Q179 Q180  DFXTP_2_10X
X10F_18 vpwr_0 VGND ff_18 Q181 Q182 Q183 Q184 Q185 Q186 Q187 Q188 Q189 Q190  DFXTP_2_10X
X10F_19 vpwr_0 VGND ff_19 Q191 Q192 Q193 Q194 Q195 Q196 Q197 Q198 Q199 Q200  DFXTP_2_10X
X10F_20 vpwr_0 VGND ff_20 Q201 Q202 Q203 Q204 Q205 Q206 Q207 Q208 Q209 Q210  DFXTP_2_10X
X10F_21 vpwr_0 VGND ff_21 Q211 Q212 Q213 Q214 Q215 Q216 Q217 Q218 Q219 Q220  DFXTP_2_10X
X10F_22 vpwr_0 VGND ff_22 Q221 Q222 Q223 Q224 Q225 Q226 Q227 Q228 Q229 Q230  DFXTP_2_10X
X10F_23 vpwr_0 VGND ff_23 Q231 Q232 Q233 Q234 Q235 Q236 Q237 Q238 Q239 Q240  DFXTP_2_10X
X10F_24 vpwr_0 VGND ff_24 Q241 Q242 Q243 Q244 Q245 Q246 Q247 Q248 Q249 Q250  DFXTP_2_10X
X10F_25 vpwr_0 VGND ff_25 Q251 Q252 Q253 Q254 Q255 Q256 Q257 Q258 Q259 Q260  DFXTP_2_10X
X10F_26 vpwr_0 VGND ff_26 Q261 Q262 Q263 Q264 Q265 Q266 Q267 Q268 Q269 Q270  DFXTP_2_10X
X10F_27 vpwr_0 VGND ff_27 Q271 Q272 Q273 Q274 Q275 Q276 Q277 Q278 Q279 Q280  DFXTP_2_10X
X10F_28 vpwr_0 VGND ff_28 Q281 Q282 Q283 Q284 Q285 Q286 Q287 Q288 Q289 Q290  DFXTP_2_10X
X10F_29 vpwr_0 VGND ff_29 Q291 Q292 Q293 Q294 Q295 Q296 Q297 Q298 Q299 Q300  DFXTP_2_10X
X10F_30 vpwr_0 VGND ff_30 Q301 Q302 Q303 Q304 Q305 Q306 Q307 Q308 Q309 Q310  DFXTP_2_10X
X10F_31 vpwr_0 VGND ff_31 Q311 Q312 Q313 Q314 Q315 Q316 Q317 Q318 Q319 Q320  DFXTP_2_10X


.lib     ../../../pdks/sky130A-1.0.227.01/libs.tech/ngspice/sky130.lib.spice ${CORNER}
.include ../../../pdks/sky130A-1.0.227.01/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include ../../dfxtp_2_10x.spice

.temp ${TEMP}
.save all
.tran 0.1n 100n

.end

magic
tech sky130A
magscale 1 2
timestamp 1633016303
<< nwell >>
rect -66 377 2754 897
<< pwell >>
rect 0 -17 2688 17
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2688 831
rect 25 729 131 751
rect 59 695 97 729
rect 25 435 131 695
rect 180 498 246 751
rect 180 464 197 498
rect 231 464 246 498
rect 19 119 126 295
rect 180 159 246 464
rect 280 729 458 751
rect 314 695 352 729
rect 386 695 424 729
rect 280 435 458 695
rect 492 498 558 751
rect 492 464 509 498
rect 543 464 558 498
rect 280 350 458 379
rect 280 316 319 350
rect 353 316 391 350
rect 425 316 458 350
rect 280 313 458 316
rect 53 85 91 119
rect 125 85 126 119
rect 19 75 126 85
rect 280 119 458 279
rect 492 159 558 464
rect 592 729 770 751
rect 626 695 664 729
rect 698 695 736 729
rect 592 435 770 695
rect 804 498 870 751
rect 804 464 821 498
rect 855 464 870 498
rect 592 350 770 379
rect 592 316 629 350
rect 663 316 701 350
rect 735 316 770 350
rect 592 313 770 316
rect 314 85 352 119
rect 386 85 424 119
rect 280 75 458 85
rect 592 119 770 279
rect 804 159 870 464
rect 904 729 1082 751
rect 938 695 976 729
rect 1010 695 1048 729
rect 904 435 1082 695
rect 1116 498 1182 751
rect 1116 464 1133 498
rect 1167 464 1182 498
rect 904 350 1082 379
rect 904 316 941 350
rect 975 316 1013 350
rect 1047 316 1082 350
rect 904 313 1082 316
rect 626 85 664 119
rect 698 85 736 119
rect 592 75 770 85
rect 904 119 1082 279
rect 1116 159 1182 464
rect 1216 729 1394 751
rect 1250 695 1288 729
rect 1322 695 1360 729
rect 1216 435 1394 695
rect 1428 498 1494 751
rect 1428 464 1445 498
rect 1479 464 1494 498
rect 1216 350 1394 379
rect 1216 316 1253 350
rect 1287 316 1325 350
rect 1359 316 1394 350
rect 1216 313 1394 316
rect 938 85 976 119
rect 1010 85 1048 119
rect 904 75 1082 85
rect 1216 119 1394 279
rect 1428 159 1494 464
rect 1528 729 1706 751
rect 1562 695 1600 729
rect 1634 695 1672 729
rect 1528 435 1706 695
rect 1740 498 1806 751
rect 1740 464 1757 498
rect 1791 464 1806 498
rect 1528 350 1706 379
rect 1528 316 1565 350
rect 1599 316 1637 350
rect 1671 316 1706 350
rect 1528 313 1706 316
rect 1250 85 1288 119
rect 1322 85 1360 119
rect 1216 75 1394 85
rect 1528 119 1706 279
rect 1740 159 1806 464
rect 1840 729 2018 751
rect 1874 695 1912 729
rect 1946 695 1984 729
rect 1840 435 2018 695
rect 2052 498 2118 751
rect 2052 464 2069 498
rect 2103 464 2118 498
rect 1840 350 2018 379
rect 1840 316 1877 350
rect 1911 316 1949 350
rect 1983 316 2018 350
rect 1840 313 2018 316
rect 1562 85 1600 119
rect 1634 85 1672 119
rect 1528 75 1706 85
rect 1840 119 2018 279
rect 2052 159 2118 464
rect 2152 729 2330 751
rect 2186 695 2224 729
rect 2258 695 2296 729
rect 2152 435 2330 695
rect 2364 498 2430 751
rect 2364 464 2381 498
rect 2415 464 2430 498
rect 2152 350 2330 379
rect 2152 316 2189 350
rect 2223 316 2261 350
rect 2295 316 2330 350
rect 2152 313 2330 316
rect 1874 85 1912 119
rect 1946 85 1984 119
rect 1840 75 2018 85
rect 2152 119 2330 279
rect 2364 159 2430 464
rect 2464 729 2587 735
rect 2464 695 2473 729
rect 2507 695 2545 729
rect 2579 695 2587 729
rect 2464 435 2587 695
rect 2186 85 2224 119
rect 2258 85 2296 119
rect 2152 75 2330 85
rect 2464 119 2587 279
rect 2464 85 2473 119
rect 2507 85 2545 119
rect 2579 85 2587 119
rect 2464 75 2587 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 25 695 59 729
rect 97 695 131 729
rect 197 464 231 498
rect 280 695 314 729
rect 352 695 386 729
rect 424 695 458 729
rect 509 464 543 498
rect 319 316 353 350
rect 391 316 425 350
rect 19 85 53 119
rect 91 85 125 119
rect 592 695 626 729
rect 664 695 698 729
rect 736 695 770 729
rect 821 464 855 498
rect 629 316 663 350
rect 701 316 735 350
rect 280 85 314 119
rect 352 85 386 119
rect 424 85 458 119
rect 904 695 938 729
rect 976 695 1010 729
rect 1048 695 1082 729
rect 1133 464 1167 498
rect 941 316 975 350
rect 1013 316 1047 350
rect 592 85 626 119
rect 664 85 698 119
rect 736 85 770 119
rect 1216 695 1250 729
rect 1288 695 1322 729
rect 1360 695 1394 729
rect 1445 464 1479 498
rect 1253 316 1287 350
rect 1325 316 1359 350
rect 904 85 938 119
rect 976 85 1010 119
rect 1048 85 1082 119
rect 1528 695 1562 729
rect 1600 695 1634 729
rect 1672 695 1706 729
rect 1757 464 1791 498
rect 1565 316 1599 350
rect 1637 316 1671 350
rect 1216 85 1250 119
rect 1288 85 1322 119
rect 1360 85 1394 119
rect 1840 695 1874 729
rect 1912 695 1946 729
rect 1984 695 2018 729
rect 2069 464 2103 498
rect 1877 316 1911 350
rect 1949 316 1983 350
rect 1528 85 1562 119
rect 1600 85 1634 119
rect 1672 85 1706 119
rect 2152 695 2186 729
rect 2224 695 2258 729
rect 2296 695 2330 729
rect 2381 464 2415 498
rect 2189 316 2223 350
rect 2261 316 2295 350
rect 1840 85 1874 119
rect 1912 85 1946 119
rect 1984 85 2018 119
rect 2473 695 2507 729
rect 2545 695 2579 729
rect 2152 85 2186 119
rect 2224 85 2258 119
rect 2296 85 2330 119
rect 2473 85 2507 119
rect 2545 85 2579 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 831 2688 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2688 831
rect 0 791 2688 797
rect 0 729 2688 763
rect 0 695 25 729
rect 59 695 97 729
rect 131 695 280 729
rect 314 695 352 729
rect 386 695 424 729
rect 458 695 592 729
rect 626 695 664 729
rect 698 695 736 729
rect 770 695 904 729
rect 938 695 976 729
rect 1010 695 1048 729
rect 1082 695 1216 729
rect 1250 695 1288 729
rect 1322 695 1360 729
rect 1394 695 1528 729
rect 1562 695 1600 729
rect 1634 695 1672 729
rect 1706 695 1840 729
rect 1874 695 1912 729
rect 1946 695 1984 729
rect 2018 695 2152 729
rect 2186 695 2224 729
rect 2258 695 2296 729
rect 2330 695 2473 729
rect 2507 695 2545 729
rect 2579 695 2688 729
rect 0 689 2688 695
rect 185 498 243 504
rect 497 498 555 504
rect 809 498 867 504
rect 1121 498 1179 504
rect 1433 498 1491 504
rect 1745 498 1803 504
rect 2057 498 2115 504
rect 2369 498 2427 504
rect 185 464 197 498
rect 231 464 509 498
rect 543 464 821 498
rect 855 464 1133 498
rect 1167 464 1445 498
rect 1479 464 1757 498
rect 1791 464 2069 498
rect 2103 464 2381 498
rect 2415 464 2427 498
rect 185 458 243 464
rect 497 458 555 464
rect 809 458 867 464
rect 1121 458 1179 464
rect 1433 458 1491 464
rect 1745 458 1803 464
rect 2057 458 2115 464
rect 2369 458 2427 464
rect 307 350 437 356
rect 617 350 747 356
rect 929 350 1059 356
rect 1241 350 1371 356
rect 1553 350 1683 356
rect 1865 350 1995 356
rect 2177 350 2307 356
rect 307 316 319 350
rect 353 316 391 350
rect 425 316 629 350
rect 663 316 701 350
rect 735 316 941 350
rect 975 316 1013 350
rect 1047 316 1253 350
rect 1287 316 1325 350
rect 1359 316 1565 350
rect 1599 316 1637 350
rect 1671 316 1877 350
rect 1911 316 1949 350
rect 1983 316 2189 350
rect 2223 316 2261 350
rect 2295 316 2307 350
rect 307 310 437 316
rect 617 310 747 316
rect 929 310 1059 316
rect 1241 310 1371 316
rect 1553 310 1683 316
rect 1865 310 1995 316
rect 2177 310 2307 316
rect 0 119 2688 125
rect 0 85 19 119
rect 53 85 91 119
rect 125 85 280 119
rect 314 85 352 119
rect 386 85 424 119
rect 458 85 592 119
rect 626 85 664 119
rect 698 85 736 119
rect 770 85 904 119
rect 938 85 976 119
rect 1010 85 1048 119
rect 1082 85 1216 119
rect 1250 85 1288 119
rect 1322 85 1360 119
rect 1394 85 1528 119
rect 1562 85 1600 119
rect 1634 85 1672 119
rect 1706 85 1840 119
rect 1874 85 1912 119
rect 1946 85 1984 119
rect 2018 85 2152 119
rect 2186 85 2224 119
rect 2258 85 2296 119
rect 2330 85 2473 119
rect 2507 85 2545 119
rect 2579 85 2688 119
rect 0 51 2688 85
rect 0 17 2688 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -23 2688 -17
<< labels >>
rlabel metal1 s 2177 350 2307 356 6 A
port 1 nsew signal input
rlabel metal1 s 2177 310 2307 316 6 A
port 1 nsew signal input
rlabel metal1 s 1865 350 1995 356 6 A
port 1 nsew signal input
rlabel metal1 s 1865 310 1995 316 6 A
port 1 nsew signal input
rlabel metal1 s 1553 350 1683 356 6 A
port 1 nsew signal input
rlabel metal1 s 1553 310 1683 316 6 A
port 1 nsew signal input
rlabel metal1 s 1241 350 1371 356 6 A
port 1 nsew signal input
rlabel metal1 s 1241 310 1371 316 6 A
port 1 nsew signal input
rlabel metal1 s 929 350 1059 356 6 A
port 1 nsew signal input
rlabel metal1 s 929 310 1059 316 6 A
port 1 nsew signal input
rlabel metal1 s 617 350 747 356 6 A
port 1 nsew signal input
rlabel metal1 s 617 310 747 316 6 A
port 1 nsew signal input
rlabel metal1 s 307 350 437 356 6 A
port 1 nsew signal input
rlabel metal1 s 307 316 2307 350 6 A
port 1 nsew signal input
rlabel metal1 s 307 310 437 316 6 A
port 1 nsew signal input
rlabel metal1 s 2369 498 2427 504 6 Y
port 6 nsew signal output
rlabel metal1 s 2369 458 2427 464 6 Y
port 6 nsew signal output
rlabel metal1 s 2057 498 2115 504 6 Y
port 6 nsew signal output
rlabel metal1 s 2057 458 2115 464 6 Y
port 6 nsew signal output
rlabel metal1 s 1745 498 1803 504 6 Y
port 6 nsew signal output
rlabel metal1 s 1745 458 1803 464 6 Y
port 6 nsew signal output
rlabel metal1 s 1433 498 1491 504 6 Y
port 6 nsew signal output
rlabel metal1 s 1433 458 1491 464 6 Y
port 6 nsew signal output
rlabel metal1 s 1121 498 1179 504 6 Y
port 6 nsew signal output
rlabel metal1 s 1121 458 1179 464 6 Y
port 6 nsew signal output
rlabel metal1 s 809 498 867 504 6 Y
port 6 nsew signal output
rlabel metal1 s 809 458 867 464 6 Y
port 6 nsew signal output
rlabel metal1 s 497 498 555 504 6 Y
port 6 nsew signal output
rlabel metal1 s 497 458 555 464 6 Y
port 6 nsew signal output
rlabel metal1 s 185 498 243 504 6 Y
port 6 nsew signal output
rlabel metal1 s 185 464 2427 498 6 Y
port 6 nsew signal output
rlabel metal1 s 185 458 243 464 6 Y
port 6 nsew signal output
rlabel metal1 s 0 51 2688 125 6 VGND
port 2 nsew ground bidirectional
rlabel pwell s 0 -17 2688 17 8 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 2688 23 8 VNB
port 3 nsew ground bidirectional
rlabel nwell s -66 377 2754 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 791 2688 837 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 2688 763 6 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 2688 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 78564
string GDS_START 48924
<< end >>

* NGSPICE file created from sky130_ef_sc_hd__fill_8.ext - technology: sky130A

.subckt sky130_ef_sc_hd__fill_8 VGND VPWR VPB VNB
C0 a_31_305# VPWR 0.14fF
C1 a_31_39# VGND 0.14fF
.ends


magic
tech sky130A
magscale 1 2
timestamp 1633016078
<< obsli1 >>
rect 34 2492 2158 2558
rect 34 100 100 2492
rect 260 2266 1932 2332
rect 260 326 326 2266
rect 662 1864 1530 1930
rect 662 728 728 1864
rect 893 893 1299 1699
rect 1464 728 1530 1864
rect 662 662 1530 728
rect 1866 326 1932 2266
rect 260 260 1932 326
rect 2092 100 2158 2492
rect 34 34 2158 100
<< obsm1 >>
rect 38 2496 2154 2554
rect 38 96 96 2496
rect 264 2270 1928 2328
rect 264 322 322 2270
rect 666 1868 1526 1926
rect 666 724 724 1868
rect 923 943 1269 1649
rect 1468 724 1526 1868
rect 666 666 1526 724
rect 1870 322 1928 2270
rect 264 264 1928 322
rect 2096 96 2154 2496
rect 38 38 2154 96
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 26 26 2166 2566
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 8734936
string GDS_START 8682124
<< end >>

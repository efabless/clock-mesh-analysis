magic
tech sky130A
magscale 1 2
timestamp 1633016303
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 0 -17 768 17
<< locali >>
rect 185 435 257 691
rect 25 301 167 367
rect 217 196 257 435
rect 293 301 359 350
rect 409 301 551 350
rect 588 301 743 350
rect 341 196 391 265
rect 217 162 391 196
rect 341 99 391 162
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 29 727 391 761
rect 29 435 95 727
rect 18 113 136 265
rect 341 420 391 727
rect 427 735 617 751
rect 427 701 433 735
rect 467 701 505 735
rect 539 701 577 735
rect 611 701 617 735
rect 427 456 617 701
rect 653 420 719 751
rect 341 386 719 420
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 136 113
rect 427 113 750 265
rect 18 73 136 79
rect 461 79 499 113
rect 533 79 571 113
rect 605 79 643 113
rect 677 79 715 113
rect 749 79 750 113
rect 427 73 750 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 433 701 467 735
rect 505 701 539 735
rect 577 701 611 735
rect 24 79 58 113
rect 96 79 130 113
rect 427 79 461 113
rect 499 79 533 113
rect 571 79 605 113
rect 643 79 677 113
rect 715 79 749 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 735 768 763
rect 0 701 433 735
rect 467 701 505 735
rect 539 701 577 735
rect 611 701 768 735
rect 0 689 768 701
rect 0 113 768 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 427 113
rect 461 79 499 113
rect 533 79 571 113
rect 605 79 643 113
rect 677 79 715 113
rect 749 79 768 113
rect 0 51 768 79
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel locali s 409 301 551 350 6 A1
port 1 nsew signal input
rlabel locali s 588 301 743 350 6 A2
port 2 nsew signal input
rlabel locali s 293 301 359 350 6 B1
port 3 nsew signal input
rlabel locali s 25 301 167 367 6 B2
port 4 nsew signal input
rlabel locali s 341 196 391 265 6 Y
port 9 nsew signal output
rlabel locali s 341 99 391 162 6 Y
port 9 nsew signal output
rlabel locali s 217 196 257 435 6 Y
port 9 nsew signal output
rlabel locali s 217 162 391 196 6 Y
port 9 nsew signal output
rlabel locali s 185 435 257 691 6 Y
port 9 nsew signal output
rlabel metal1 s 0 51 768 125 6 VGND
port 5 nsew ground bidirectional
rlabel pwell s 0 -17 768 17 8 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 -23 768 23 8 VNB
port 6 nsew ground bidirectional
rlabel nwell s -66 377 834 897 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 791 768 837 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 689 768 763 6 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 768 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 789130
string GDS_START 778648
<< end >>

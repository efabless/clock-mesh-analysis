magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -2107 -4091 13331 3119
<< dnwell >>
rect 26 30 11991 1672
<< nwell >>
rect -54 1466 12071 1752
rect -54 236 232 1466
rect 1839 236 2075 1466
rect 6817 236 7053 1466
rect -54 -50 12071 236
rect 5550 -1087 7628 -1086
rect 5550 -2111 8043 -1087
<< pwell >>
rect 331 296 1735 1380
rect 2166 296 6726 1406
rect 7170 296 11744 1406
<< mvnmos >>
rect 558 1087 1558 1187
rect 558 931 1558 1031
rect 558 645 1558 745
rect 558 489 1558 589
rect 2393 1113 4393 1213
rect 4499 1113 6499 1213
rect 2393 957 4393 1057
rect 4499 957 6499 1057
rect 2393 801 4393 901
rect 4499 801 6499 901
rect 2393 645 4393 745
rect 4499 645 6499 745
rect 2393 489 4393 589
rect 4499 489 6499 589
rect 7412 1113 9412 1213
rect 9518 1113 11518 1213
rect 7412 957 9412 1057
rect 9518 957 11518 1057
rect 7412 801 9412 901
rect 9518 801 11518 901
rect 7412 645 9412 745
rect 9518 645 11518 745
rect 7412 489 9412 589
rect 9518 489 11518 589
<< mvpmos >>
rect 5816 -1415 7816 -1315
rect 5816 -1571 7816 -1471
rect 5816 -1727 7816 -1627
rect 5816 -1883 7816 -1783
<< mvndiff >>
rect 558 1232 1558 1240
rect 558 1198 570 1232
rect 604 1198 638 1232
rect 672 1198 706 1232
rect 740 1198 774 1232
rect 808 1198 842 1232
rect 876 1198 910 1232
rect 944 1198 978 1232
rect 1012 1198 1046 1232
rect 1080 1198 1114 1232
rect 1148 1198 1182 1232
rect 1216 1198 1250 1232
rect 1284 1198 1318 1232
rect 1352 1198 1386 1232
rect 1420 1198 1454 1232
rect 1488 1198 1558 1232
rect 558 1187 1558 1198
rect 558 1076 1558 1087
rect 558 1042 570 1076
rect 604 1042 638 1076
rect 672 1042 706 1076
rect 740 1042 774 1076
rect 808 1042 842 1076
rect 876 1042 910 1076
rect 944 1042 978 1076
rect 1012 1042 1046 1076
rect 1080 1042 1114 1076
rect 1148 1042 1182 1076
rect 1216 1042 1250 1076
rect 1284 1042 1318 1076
rect 1352 1042 1386 1076
rect 1420 1042 1454 1076
rect 1488 1042 1558 1076
rect 558 1031 1558 1042
rect 558 920 1558 931
rect 558 886 570 920
rect 604 886 638 920
rect 672 886 706 920
rect 740 886 774 920
rect 808 886 842 920
rect 876 886 910 920
rect 944 886 978 920
rect 1012 886 1046 920
rect 1080 886 1114 920
rect 1148 886 1182 920
rect 1216 886 1250 920
rect 1284 886 1318 920
rect 1352 886 1386 920
rect 1420 886 1454 920
rect 1488 886 1558 920
rect 558 878 1558 886
rect 558 790 1558 798
rect 558 756 570 790
rect 604 756 638 790
rect 672 756 706 790
rect 740 756 774 790
rect 808 756 842 790
rect 876 756 910 790
rect 944 756 978 790
rect 1012 756 1046 790
rect 1080 756 1114 790
rect 1148 756 1182 790
rect 1216 756 1250 790
rect 1284 756 1318 790
rect 1352 756 1386 790
rect 1420 756 1454 790
rect 1488 756 1558 790
rect 558 745 1558 756
rect 558 634 1558 645
rect 558 600 570 634
rect 604 600 638 634
rect 672 600 706 634
rect 740 600 774 634
rect 808 600 842 634
rect 876 600 910 634
rect 944 600 978 634
rect 1012 600 1046 634
rect 1080 600 1114 634
rect 1148 600 1182 634
rect 1216 600 1250 634
rect 1284 600 1318 634
rect 1352 600 1386 634
rect 1420 600 1454 634
rect 1488 600 1558 634
rect 558 589 1558 600
rect 558 478 1558 489
rect 558 444 570 478
rect 604 444 638 478
rect 672 444 706 478
rect 740 444 774 478
rect 808 444 842 478
rect 876 444 910 478
rect 944 444 978 478
rect 1012 444 1046 478
rect 1080 444 1114 478
rect 1148 444 1182 478
rect 1216 444 1250 478
rect 1284 444 1318 478
rect 1352 444 1386 478
rect 1420 444 1454 478
rect 1488 444 1558 478
rect 558 436 1558 444
rect 2393 1258 4393 1266
rect 2393 1224 2405 1258
rect 2439 1224 2473 1258
rect 2507 1224 2541 1258
rect 2575 1224 2609 1258
rect 2643 1224 2677 1258
rect 2711 1224 2745 1258
rect 2779 1224 2813 1258
rect 2847 1224 2881 1258
rect 2915 1224 2949 1258
rect 2983 1224 3017 1258
rect 3051 1224 3085 1258
rect 3119 1224 3153 1258
rect 3187 1224 3221 1258
rect 3255 1224 3289 1258
rect 3323 1224 3357 1258
rect 3391 1224 3425 1258
rect 3459 1224 3493 1258
rect 3527 1224 3561 1258
rect 3595 1224 3629 1258
rect 3663 1224 3697 1258
rect 3731 1224 3765 1258
rect 3799 1224 3833 1258
rect 3867 1224 3901 1258
rect 3935 1224 3969 1258
rect 4003 1224 4037 1258
rect 4071 1224 4105 1258
rect 4139 1224 4173 1258
rect 4207 1224 4241 1258
rect 4275 1224 4309 1258
rect 4343 1224 4393 1258
rect 2393 1213 4393 1224
rect 4499 1258 6499 1266
rect 4499 1224 4549 1258
rect 4583 1224 4617 1258
rect 4651 1224 4685 1258
rect 4719 1224 4753 1258
rect 4787 1224 4821 1258
rect 4855 1224 4889 1258
rect 4923 1224 4957 1258
rect 4991 1224 5025 1258
rect 5059 1224 5093 1258
rect 5127 1224 5161 1258
rect 5195 1224 5229 1258
rect 5263 1224 5297 1258
rect 5331 1224 5365 1258
rect 5399 1224 5433 1258
rect 5467 1224 5501 1258
rect 5535 1224 5569 1258
rect 5603 1224 5637 1258
rect 5671 1224 5705 1258
rect 5739 1224 5773 1258
rect 5807 1224 5841 1258
rect 5875 1224 5909 1258
rect 5943 1224 5977 1258
rect 6011 1224 6045 1258
rect 6079 1224 6113 1258
rect 6147 1224 6181 1258
rect 6215 1224 6249 1258
rect 6283 1224 6317 1258
rect 6351 1224 6385 1258
rect 6419 1224 6453 1258
rect 6487 1224 6499 1258
rect 4499 1213 6499 1224
rect 2393 1102 4393 1113
rect 2393 1068 2405 1102
rect 2439 1068 2473 1102
rect 2507 1068 2541 1102
rect 2575 1068 2609 1102
rect 2643 1068 2677 1102
rect 2711 1068 2745 1102
rect 2779 1068 2813 1102
rect 2847 1068 2881 1102
rect 2915 1068 2949 1102
rect 2983 1068 3017 1102
rect 3051 1068 3085 1102
rect 3119 1068 3153 1102
rect 3187 1068 3221 1102
rect 3255 1068 3289 1102
rect 3323 1068 3357 1102
rect 3391 1068 3425 1102
rect 3459 1068 3493 1102
rect 3527 1068 3561 1102
rect 3595 1068 3629 1102
rect 3663 1068 3697 1102
rect 3731 1068 3765 1102
rect 3799 1068 3833 1102
rect 3867 1068 3901 1102
rect 3935 1068 3969 1102
rect 4003 1068 4037 1102
rect 4071 1068 4105 1102
rect 4139 1068 4173 1102
rect 4207 1068 4241 1102
rect 4275 1068 4309 1102
rect 4343 1068 4393 1102
rect 2393 1057 4393 1068
rect 4499 1102 6499 1113
rect 4499 1068 4549 1102
rect 4583 1068 4617 1102
rect 4651 1068 4685 1102
rect 4719 1068 4753 1102
rect 4787 1068 4821 1102
rect 4855 1068 4889 1102
rect 4923 1068 4957 1102
rect 4991 1068 5025 1102
rect 5059 1068 5093 1102
rect 5127 1068 5161 1102
rect 5195 1068 5229 1102
rect 5263 1068 5297 1102
rect 5331 1068 5365 1102
rect 5399 1068 5433 1102
rect 5467 1068 5501 1102
rect 5535 1068 5569 1102
rect 5603 1068 5637 1102
rect 5671 1068 5705 1102
rect 5739 1068 5773 1102
rect 5807 1068 5841 1102
rect 5875 1068 5909 1102
rect 5943 1068 5977 1102
rect 6011 1068 6045 1102
rect 6079 1068 6113 1102
rect 6147 1068 6181 1102
rect 6215 1068 6249 1102
rect 6283 1068 6317 1102
rect 6351 1068 6385 1102
rect 6419 1068 6453 1102
rect 6487 1068 6499 1102
rect 4499 1057 6499 1068
rect 2393 946 4393 957
rect 2393 912 2405 946
rect 2439 912 2473 946
rect 2507 912 2541 946
rect 2575 912 2609 946
rect 2643 912 2677 946
rect 2711 912 2745 946
rect 2779 912 2813 946
rect 2847 912 2881 946
rect 2915 912 2949 946
rect 2983 912 3017 946
rect 3051 912 3085 946
rect 3119 912 3153 946
rect 3187 912 3221 946
rect 3255 912 3289 946
rect 3323 912 3357 946
rect 3391 912 3425 946
rect 3459 912 3493 946
rect 3527 912 3561 946
rect 3595 912 3629 946
rect 3663 912 3697 946
rect 3731 912 3765 946
rect 3799 912 3833 946
rect 3867 912 3901 946
rect 3935 912 3969 946
rect 4003 912 4037 946
rect 4071 912 4105 946
rect 4139 912 4173 946
rect 4207 912 4241 946
rect 4275 912 4309 946
rect 4343 912 4393 946
rect 2393 901 4393 912
rect 4499 946 6499 957
rect 4499 912 4549 946
rect 4583 912 4617 946
rect 4651 912 4685 946
rect 4719 912 4753 946
rect 4787 912 4821 946
rect 4855 912 4889 946
rect 4923 912 4957 946
rect 4991 912 5025 946
rect 5059 912 5093 946
rect 5127 912 5161 946
rect 5195 912 5229 946
rect 5263 912 5297 946
rect 5331 912 5365 946
rect 5399 912 5433 946
rect 5467 912 5501 946
rect 5535 912 5569 946
rect 5603 912 5637 946
rect 5671 912 5705 946
rect 5739 912 5773 946
rect 5807 912 5841 946
rect 5875 912 5909 946
rect 5943 912 5977 946
rect 6011 912 6045 946
rect 6079 912 6113 946
rect 6147 912 6181 946
rect 6215 912 6249 946
rect 6283 912 6317 946
rect 6351 912 6385 946
rect 6419 912 6453 946
rect 6487 912 6499 946
rect 4499 901 6499 912
rect 2393 790 4393 801
rect 2393 756 2405 790
rect 2439 756 2473 790
rect 2507 756 2541 790
rect 2575 756 2609 790
rect 2643 756 2677 790
rect 2711 756 2745 790
rect 2779 756 2813 790
rect 2847 756 2881 790
rect 2915 756 2949 790
rect 2983 756 3017 790
rect 3051 756 3085 790
rect 3119 756 3153 790
rect 3187 756 3221 790
rect 3255 756 3289 790
rect 3323 756 3357 790
rect 3391 756 3425 790
rect 3459 756 3493 790
rect 3527 756 3561 790
rect 3595 756 3629 790
rect 3663 756 3697 790
rect 3731 756 3765 790
rect 3799 756 3833 790
rect 3867 756 3901 790
rect 3935 756 3969 790
rect 4003 756 4037 790
rect 4071 756 4105 790
rect 4139 756 4173 790
rect 4207 756 4241 790
rect 4275 756 4309 790
rect 4343 756 4393 790
rect 2393 745 4393 756
rect 4499 790 6499 801
rect 4499 756 4549 790
rect 4583 756 4617 790
rect 4651 756 4685 790
rect 4719 756 4753 790
rect 4787 756 4821 790
rect 4855 756 4889 790
rect 4923 756 4957 790
rect 4991 756 5025 790
rect 5059 756 5093 790
rect 5127 756 5161 790
rect 5195 756 5229 790
rect 5263 756 5297 790
rect 5331 756 5365 790
rect 5399 756 5433 790
rect 5467 756 5501 790
rect 5535 756 5569 790
rect 5603 756 5637 790
rect 5671 756 5705 790
rect 5739 756 5773 790
rect 5807 756 5841 790
rect 5875 756 5909 790
rect 5943 756 5977 790
rect 6011 756 6045 790
rect 6079 756 6113 790
rect 6147 756 6181 790
rect 6215 756 6249 790
rect 6283 756 6317 790
rect 6351 756 6385 790
rect 6419 756 6453 790
rect 6487 756 6499 790
rect 4499 745 6499 756
rect 2393 634 4393 645
rect 2393 600 2405 634
rect 2439 600 2473 634
rect 2507 600 2541 634
rect 2575 600 2609 634
rect 2643 600 2677 634
rect 2711 600 2745 634
rect 2779 600 2813 634
rect 2847 600 2881 634
rect 2915 600 2949 634
rect 2983 600 3017 634
rect 3051 600 3085 634
rect 3119 600 3153 634
rect 3187 600 3221 634
rect 3255 600 3289 634
rect 3323 600 3357 634
rect 3391 600 3425 634
rect 3459 600 3493 634
rect 3527 600 3561 634
rect 3595 600 3629 634
rect 3663 600 3697 634
rect 3731 600 3765 634
rect 3799 600 3833 634
rect 3867 600 3901 634
rect 3935 600 3969 634
rect 4003 600 4037 634
rect 4071 600 4105 634
rect 4139 600 4173 634
rect 4207 600 4241 634
rect 4275 600 4309 634
rect 4343 600 4393 634
rect 2393 589 4393 600
rect 4499 634 6499 645
rect 4499 600 4549 634
rect 4583 600 4617 634
rect 4651 600 4685 634
rect 4719 600 4753 634
rect 4787 600 4821 634
rect 4855 600 4889 634
rect 4923 600 4957 634
rect 4991 600 5025 634
rect 5059 600 5093 634
rect 5127 600 5161 634
rect 5195 600 5229 634
rect 5263 600 5297 634
rect 5331 600 5365 634
rect 5399 600 5433 634
rect 5467 600 5501 634
rect 5535 600 5569 634
rect 5603 600 5637 634
rect 5671 600 5705 634
rect 5739 600 5773 634
rect 5807 600 5841 634
rect 5875 600 5909 634
rect 5943 600 5977 634
rect 6011 600 6045 634
rect 6079 600 6113 634
rect 6147 600 6181 634
rect 6215 600 6249 634
rect 6283 600 6317 634
rect 6351 600 6385 634
rect 6419 600 6453 634
rect 6487 600 6499 634
rect 4499 589 6499 600
rect 2393 478 4393 489
rect 2393 444 2405 478
rect 2439 444 2473 478
rect 2507 444 2541 478
rect 2575 444 2609 478
rect 2643 444 2677 478
rect 2711 444 2745 478
rect 2779 444 2813 478
rect 2847 444 2881 478
rect 2915 444 2949 478
rect 2983 444 3017 478
rect 3051 444 3085 478
rect 3119 444 3153 478
rect 3187 444 3221 478
rect 3255 444 3289 478
rect 3323 444 3357 478
rect 3391 444 3425 478
rect 3459 444 3493 478
rect 3527 444 3561 478
rect 3595 444 3629 478
rect 3663 444 3697 478
rect 3731 444 3765 478
rect 3799 444 3833 478
rect 3867 444 3901 478
rect 3935 444 3969 478
rect 4003 444 4037 478
rect 4071 444 4105 478
rect 4139 444 4173 478
rect 4207 444 4241 478
rect 4275 444 4309 478
rect 4343 444 4393 478
rect 2393 436 4393 444
rect 4499 478 6499 489
rect 4499 444 4549 478
rect 4583 444 4617 478
rect 4651 444 4685 478
rect 4719 444 4753 478
rect 4787 444 4821 478
rect 4855 444 4889 478
rect 4923 444 4957 478
rect 4991 444 5025 478
rect 5059 444 5093 478
rect 5127 444 5161 478
rect 5195 444 5229 478
rect 5263 444 5297 478
rect 5331 444 5365 478
rect 5399 444 5433 478
rect 5467 444 5501 478
rect 5535 444 5569 478
rect 5603 444 5637 478
rect 5671 444 5705 478
rect 5739 444 5773 478
rect 5807 444 5841 478
rect 5875 444 5909 478
rect 5943 444 5977 478
rect 6011 444 6045 478
rect 6079 444 6113 478
rect 6147 444 6181 478
rect 6215 444 6249 478
rect 6283 444 6317 478
rect 6351 444 6385 478
rect 6419 444 6453 478
rect 6487 444 6499 478
rect 4499 436 6499 444
rect 7412 1258 9412 1266
rect 7412 1224 7462 1258
rect 7496 1224 7530 1258
rect 7564 1224 7598 1258
rect 7632 1224 7666 1258
rect 7700 1224 7734 1258
rect 7768 1224 7802 1258
rect 7836 1224 7870 1258
rect 7904 1224 7938 1258
rect 7972 1224 8006 1258
rect 8040 1224 8074 1258
rect 8108 1224 8142 1258
rect 8176 1224 8210 1258
rect 8244 1224 8278 1258
rect 8312 1224 8346 1258
rect 8380 1224 8414 1258
rect 8448 1224 8482 1258
rect 8516 1224 8550 1258
rect 8584 1224 8618 1258
rect 8652 1224 8686 1258
rect 8720 1224 8754 1258
rect 8788 1224 8822 1258
rect 8856 1224 8890 1258
rect 8924 1224 8958 1258
rect 8992 1224 9026 1258
rect 9060 1224 9094 1258
rect 9128 1224 9162 1258
rect 9196 1224 9230 1258
rect 9264 1224 9298 1258
rect 9332 1224 9366 1258
rect 9400 1224 9412 1258
rect 7412 1213 9412 1224
rect 9518 1258 11518 1266
rect 9518 1224 9568 1258
rect 9602 1224 9636 1258
rect 9670 1224 9704 1258
rect 9738 1224 9772 1258
rect 9806 1224 9840 1258
rect 9874 1224 9908 1258
rect 9942 1224 9976 1258
rect 10010 1224 10044 1258
rect 10078 1224 10112 1258
rect 10146 1224 10180 1258
rect 10214 1224 10248 1258
rect 10282 1224 10316 1258
rect 10350 1224 10384 1258
rect 10418 1224 10452 1258
rect 10486 1224 10520 1258
rect 10554 1224 10588 1258
rect 10622 1224 10656 1258
rect 10690 1224 10724 1258
rect 10758 1224 10792 1258
rect 10826 1224 10860 1258
rect 10894 1224 10928 1258
rect 10962 1224 10996 1258
rect 11030 1224 11064 1258
rect 11098 1224 11132 1258
rect 11166 1224 11200 1258
rect 11234 1224 11268 1258
rect 11302 1224 11336 1258
rect 11370 1224 11404 1258
rect 11438 1224 11472 1258
rect 11506 1224 11518 1258
rect 9518 1213 11518 1224
rect 7412 1102 9412 1113
rect 7412 1068 7462 1102
rect 7496 1068 7530 1102
rect 7564 1068 7598 1102
rect 7632 1068 7666 1102
rect 7700 1068 7734 1102
rect 7768 1068 7802 1102
rect 7836 1068 7870 1102
rect 7904 1068 7938 1102
rect 7972 1068 8006 1102
rect 8040 1068 8074 1102
rect 8108 1068 8142 1102
rect 8176 1068 8210 1102
rect 8244 1068 8278 1102
rect 8312 1068 8346 1102
rect 8380 1068 8414 1102
rect 8448 1068 8482 1102
rect 8516 1068 8550 1102
rect 8584 1068 8618 1102
rect 8652 1068 8686 1102
rect 8720 1068 8754 1102
rect 8788 1068 8822 1102
rect 8856 1068 8890 1102
rect 8924 1068 8958 1102
rect 8992 1068 9026 1102
rect 9060 1068 9094 1102
rect 9128 1068 9162 1102
rect 9196 1068 9230 1102
rect 9264 1068 9298 1102
rect 9332 1068 9366 1102
rect 9400 1068 9412 1102
rect 7412 1057 9412 1068
rect 9518 1102 11518 1113
rect 9518 1068 9568 1102
rect 9602 1068 9636 1102
rect 9670 1068 9704 1102
rect 9738 1068 9772 1102
rect 9806 1068 9840 1102
rect 9874 1068 9908 1102
rect 9942 1068 9976 1102
rect 10010 1068 10044 1102
rect 10078 1068 10112 1102
rect 10146 1068 10180 1102
rect 10214 1068 10248 1102
rect 10282 1068 10316 1102
rect 10350 1068 10384 1102
rect 10418 1068 10452 1102
rect 10486 1068 10520 1102
rect 10554 1068 10588 1102
rect 10622 1068 10656 1102
rect 10690 1068 10724 1102
rect 10758 1068 10792 1102
rect 10826 1068 10860 1102
rect 10894 1068 10928 1102
rect 10962 1068 10996 1102
rect 11030 1068 11064 1102
rect 11098 1068 11132 1102
rect 11166 1068 11200 1102
rect 11234 1068 11268 1102
rect 11302 1068 11336 1102
rect 11370 1068 11404 1102
rect 11438 1068 11472 1102
rect 11506 1068 11518 1102
rect 9518 1057 11518 1068
rect 7412 946 9412 957
rect 7412 912 7462 946
rect 7496 912 7530 946
rect 7564 912 7598 946
rect 7632 912 7666 946
rect 7700 912 7734 946
rect 7768 912 7802 946
rect 7836 912 7870 946
rect 7904 912 7938 946
rect 7972 912 8006 946
rect 8040 912 8074 946
rect 8108 912 8142 946
rect 8176 912 8210 946
rect 8244 912 8278 946
rect 8312 912 8346 946
rect 8380 912 8414 946
rect 8448 912 8482 946
rect 8516 912 8550 946
rect 8584 912 8618 946
rect 8652 912 8686 946
rect 8720 912 8754 946
rect 8788 912 8822 946
rect 8856 912 8890 946
rect 8924 912 8958 946
rect 8992 912 9026 946
rect 9060 912 9094 946
rect 9128 912 9162 946
rect 9196 912 9230 946
rect 9264 912 9298 946
rect 9332 912 9366 946
rect 9400 912 9412 946
rect 7412 901 9412 912
rect 9518 946 11518 957
rect 9518 912 9568 946
rect 9602 912 9636 946
rect 9670 912 9704 946
rect 9738 912 9772 946
rect 9806 912 9840 946
rect 9874 912 9908 946
rect 9942 912 9976 946
rect 10010 912 10044 946
rect 10078 912 10112 946
rect 10146 912 10180 946
rect 10214 912 10248 946
rect 10282 912 10316 946
rect 10350 912 10384 946
rect 10418 912 10452 946
rect 10486 912 10520 946
rect 10554 912 10588 946
rect 10622 912 10656 946
rect 10690 912 10724 946
rect 10758 912 10792 946
rect 10826 912 10860 946
rect 10894 912 10928 946
rect 10962 912 10996 946
rect 11030 912 11064 946
rect 11098 912 11132 946
rect 11166 912 11200 946
rect 11234 912 11268 946
rect 11302 912 11336 946
rect 11370 912 11404 946
rect 11438 912 11472 946
rect 11506 912 11518 946
rect 9518 901 11518 912
rect 7412 790 9412 801
rect 7412 756 7462 790
rect 7496 756 7530 790
rect 7564 756 7598 790
rect 7632 756 7666 790
rect 7700 756 7734 790
rect 7768 756 7802 790
rect 7836 756 7870 790
rect 7904 756 7938 790
rect 7972 756 8006 790
rect 8040 756 8074 790
rect 8108 756 8142 790
rect 8176 756 8210 790
rect 8244 756 8278 790
rect 8312 756 8346 790
rect 8380 756 8414 790
rect 8448 756 8482 790
rect 8516 756 8550 790
rect 8584 756 8618 790
rect 8652 756 8686 790
rect 8720 756 8754 790
rect 8788 756 8822 790
rect 8856 756 8890 790
rect 8924 756 8958 790
rect 8992 756 9026 790
rect 9060 756 9094 790
rect 9128 756 9162 790
rect 9196 756 9230 790
rect 9264 756 9298 790
rect 9332 756 9366 790
rect 9400 756 9412 790
rect 7412 745 9412 756
rect 9518 790 11518 801
rect 9518 756 9568 790
rect 9602 756 9636 790
rect 9670 756 9704 790
rect 9738 756 9772 790
rect 9806 756 9840 790
rect 9874 756 9908 790
rect 9942 756 9976 790
rect 10010 756 10044 790
rect 10078 756 10112 790
rect 10146 756 10180 790
rect 10214 756 10248 790
rect 10282 756 10316 790
rect 10350 756 10384 790
rect 10418 756 10452 790
rect 10486 756 10520 790
rect 10554 756 10588 790
rect 10622 756 10656 790
rect 10690 756 10724 790
rect 10758 756 10792 790
rect 10826 756 10860 790
rect 10894 756 10928 790
rect 10962 756 10996 790
rect 11030 756 11064 790
rect 11098 756 11132 790
rect 11166 756 11200 790
rect 11234 756 11268 790
rect 11302 756 11336 790
rect 11370 756 11404 790
rect 11438 756 11472 790
rect 11506 756 11518 790
rect 9518 745 11518 756
rect 7412 634 9412 645
rect 7412 600 7462 634
rect 7496 600 7530 634
rect 7564 600 7598 634
rect 7632 600 7666 634
rect 7700 600 7734 634
rect 7768 600 7802 634
rect 7836 600 7870 634
rect 7904 600 7938 634
rect 7972 600 8006 634
rect 8040 600 8074 634
rect 8108 600 8142 634
rect 8176 600 8210 634
rect 8244 600 8278 634
rect 8312 600 8346 634
rect 8380 600 8414 634
rect 8448 600 8482 634
rect 8516 600 8550 634
rect 8584 600 8618 634
rect 8652 600 8686 634
rect 8720 600 8754 634
rect 8788 600 8822 634
rect 8856 600 8890 634
rect 8924 600 8958 634
rect 8992 600 9026 634
rect 9060 600 9094 634
rect 9128 600 9162 634
rect 9196 600 9230 634
rect 9264 600 9298 634
rect 9332 600 9366 634
rect 9400 600 9412 634
rect 7412 589 9412 600
rect 9518 634 11518 645
rect 9518 600 9568 634
rect 9602 600 9636 634
rect 9670 600 9704 634
rect 9738 600 9772 634
rect 9806 600 9840 634
rect 9874 600 9908 634
rect 9942 600 9976 634
rect 10010 600 10044 634
rect 10078 600 10112 634
rect 10146 600 10180 634
rect 10214 600 10248 634
rect 10282 600 10316 634
rect 10350 600 10384 634
rect 10418 600 10452 634
rect 10486 600 10520 634
rect 10554 600 10588 634
rect 10622 600 10656 634
rect 10690 600 10724 634
rect 10758 600 10792 634
rect 10826 600 10860 634
rect 10894 600 10928 634
rect 10962 600 10996 634
rect 11030 600 11064 634
rect 11098 600 11132 634
rect 11166 600 11200 634
rect 11234 600 11268 634
rect 11302 600 11336 634
rect 11370 600 11404 634
rect 11438 600 11472 634
rect 11506 600 11518 634
rect 9518 589 11518 600
rect 7412 478 9412 489
rect 7412 444 7462 478
rect 7496 444 7530 478
rect 7564 444 7598 478
rect 7632 444 7666 478
rect 7700 444 7734 478
rect 7768 444 7802 478
rect 7836 444 7870 478
rect 7904 444 7938 478
rect 7972 444 8006 478
rect 8040 444 8074 478
rect 8108 444 8142 478
rect 8176 444 8210 478
rect 8244 444 8278 478
rect 8312 444 8346 478
rect 8380 444 8414 478
rect 8448 444 8482 478
rect 8516 444 8550 478
rect 8584 444 8618 478
rect 8652 444 8686 478
rect 8720 444 8754 478
rect 8788 444 8822 478
rect 8856 444 8890 478
rect 8924 444 8958 478
rect 8992 444 9026 478
rect 9060 444 9094 478
rect 9128 444 9162 478
rect 9196 444 9230 478
rect 9264 444 9298 478
rect 9332 444 9366 478
rect 9400 444 9412 478
rect 7412 436 9412 444
rect 9518 478 11518 489
rect 9518 444 9568 478
rect 9602 444 9636 478
rect 9670 444 9704 478
rect 9738 444 9772 478
rect 9806 444 9840 478
rect 9874 444 9908 478
rect 9942 444 9976 478
rect 10010 444 10044 478
rect 10078 444 10112 478
rect 10146 444 10180 478
rect 10214 444 10248 478
rect 10282 444 10316 478
rect 10350 444 10384 478
rect 10418 444 10452 478
rect 10486 444 10520 478
rect 10554 444 10588 478
rect 10622 444 10656 478
rect 10690 444 10724 478
rect 10758 444 10792 478
rect 10826 444 10860 478
rect 10894 444 10928 478
rect 10962 444 10996 478
rect 11030 444 11064 478
rect 11098 444 11132 478
rect 11166 444 11200 478
rect 11234 444 11268 478
rect 11302 444 11336 478
rect 11370 444 11404 478
rect 11438 444 11472 478
rect 11506 444 11518 478
rect 9518 436 11518 444
<< mvpdiff >>
rect 5816 -1270 7816 -1262
rect 5816 -1304 5866 -1270
rect 5900 -1304 5934 -1270
rect 5968 -1304 6002 -1270
rect 6036 -1304 6070 -1270
rect 6104 -1304 6138 -1270
rect 6172 -1304 6206 -1270
rect 6240 -1304 6274 -1270
rect 6308 -1304 6342 -1270
rect 6376 -1304 6410 -1270
rect 6444 -1304 6478 -1270
rect 6512 -1304 6546 -1270
rect 6580 -1304 6614 -1270
rect 6648 -1304 6682 -1270
rect 6716 -1304 6750 -1270
rect 6784 -1304 6818 -1270
rect 6852 -1304 6886 -1270
rect 6920 -1304 6954 -1270
rect 6988 -1304 7022 -1270
rect 7056 -1304 7090 -1270
rect 7124 -1304 7158 -1270
rect 7192 -1304 7226 -1270
rect 7260 -1304 7294 -1270
rect 7328 -1304 7362 -1270
rect 7396 -1304 7430 -1270
rect 7464 -1304 7498 -1270
rect 7532 -1304 7566 -1270
rect 7600 -1304 7634 -1270
rect 7668 -1304 7702 -1270
rect 7736 -1304 7770 -1270
rect 7804 -1304 7816 -1270
rect 5816 -1315 7816 -1304
rect 5816 -1426 7816 -1415
rect 5816 -1460 5866 -1426
rect 5900 -1460 5934 -1426
rect 5968 -1460 6002 -1426
rect 6036 -1460 6070 -1426
rect 6104 -1460 6138 -1426
rect 6172 -1460 6206 -1426
rect 6240 -1460 6274 -1426
rect 6308 -1460 6342 -1426
rect 6376 -1460 6410 -1426
rect 6444 -1460 6478 -1426
rect 6512 -1460 6546 -1426
rect 6580 -1460 6614 -1426
rect 6648 -1460 6682 -1426
rect 6716 -1460 6750 -1426
rect 6784 -1460 6818 -1426
rect 6852 -1460 6886 -1426
rect 6920 -1460 6954 -1426
rect 6988 -1460 7022 -1426
rect 7056 -1460 7090 -1426
rect 7124 -1460 7158 -1426
rect 7192 -1460 7226 -1426
rect 7260 -1460 7294 -1426
rect 7328 -1460 7362 -1426
rect 7396 -1460 7430 -1426
rect 7464 -1460 7498 -1426
rect 7532 -1460 7566 -1426
rect 7600 -1460 7634 -1426
rect 7668 -1460 7702 -1426
rect 7736 -1460 7770 -1426
rect 7804 -1460 7816 -1426
rect 5816 -1471 7816 -1460
rect 5816 -1582 7816 -1571
rect 5816 -1616 5866 -1582
rect 5900 -1616 5934 -1582
rect 5968 -1616 6002 -1582
rect 6036 -1616 6070 -1582
rect 6104 -1616 6138 -1582
rect 6172 -1616 6206 -1582
rect 6240 -1616 6274 -1582
rect 6308 -1616 6342 -1582
rect 6376 -1616 6410 -1582
rect 6444 -1616 6478 -1582
rect 6512 -1616 6546 -1582
rect 6580 -1616 6614 -1582
rect 6648 -1616 6682 -1582
rect 6716 -1616 6750 -1582
rect 6784 -1616 6818 -1582
rect 6852 -1616 6886 -1582
rect 6920 -1616 6954 -1582
rect 6988 -1616 7022 -1582
rect 7056 -1616 7090 -1582
rect 7124 -1616 7158 -1582
rect 7192 -1616 7226 -1582
rect 7260 -1616 7294 -1582
rect 7328 -1616 7362 -1582
rect 7396 -1616 7430 -1582
rect 7464 -1616 7498 -1582
rect 7532 -1616 7566 -1582
rect 7600 -1616 7634 -1582
rect 7668 -1616 7702 -1582
rect 7736 -1616 7770 -1582
rect 7804 -1616 7816 -1582
rect 5816 -1627 7816 -1616
rect 5816 -1738 7816 -1727
rect 5816 -1772 5866 -1738
rect 5900 -1772 5934 -1738
rect 5968 -1772 6002 -1738
rect 6036 -1772 6070 -1738
rect 6104 -1772 6138 -1738
rect 6172 -1772 6206 -1738
rect 6240 -1772 6274 -1738
rect 6308 -1772 6342 -1738
rect 6376 -1772 6410 -1738
rect 6444 -1772 6478 -1738
rect 6512 -1772 6546 -1738
rect 6580 -1772 6614 -1738
rect 6648 -1772 6682 -1738
rect 6716 -1772 6750 -1738
rect 6784 -1772 6818 -1738
rect 6852 -1772 6886 -1738
rect 6920 -1772 6954 -1738
rect 6988 -1772 7022 -1738
rect 7056 -1772 7090 -1738
rect 7124 -1772 7158 -1738
rect 7192 -1772 7226 -1738
rect 7260 -1772 7294 -1738
rect 7328 -1772 7362 -1738
rect 7396 -1772 7430 -1738
rect 7464 -1772 7498 -1738
rect 7532 -1772 7566 -1738
rect 7600 -1772 7634 -1738
rect 7668 -1772 7702 -1738
rect 7736 -1772 7770 -1738
rect 7804 -1772 7816 -1738
rect 5816 -1783 7816 -1772
rect 5816 -1894 7816 -1883
rect 5816 -1928 5866 -1894
rect 5900 -1928 5934 -1894
rect 5968 -1928 6002 -1894
rect 6036 -1928 6070 -1894
rect 6104 -1928 6138 -1894
rect 6172 -1928 6206 -1894
rect 6240 -1928 6274 -1894
rect 6308 -1928 6342 -1894
rect 6376 -1928 6410 -1894
rect 6444 -1928 6478 -1894
rect 6512 -1928 6546 -1894
rect 6580 -1928 6614 -1894
rect 6648 -1928 6682 -1894
rect 6716 -1928 6750 -1894
rect 6784 -1928 6818 -1894
rect 6852 -1928 6886 -1894
rect 6920 -1928 6954 -1894
rect 6988 -1928 7022 -1894
rect 7056 -1928 7090 -1894
rect 7124 -1928 7158 -1894
rect 7192 -1928 7226 -1894
rect 7260 -1928 7294 -1894
rect 7328 -1928 7362 -1894
rect 7396 -1928 7430 -1894
rect 7464 -1928 7498 -1894
rect 7532 -1928 7566 -1894
rect 7600 -1928 7634 -1894
rect 7668 -1928 7702 -1894
rect 7736 -1928 7770 -1894
rect 7804 -1928 7816 -1894
rect 5816 -1936 7816 -1928
<< mvndiffc >>
rect 570 1198 604 1232
rect 638 1198 672 1232
rect 706 1198 740 1232
rect 774 1198 808 1232
rect 842 1198 876 1232
rect 910 1198 944 1232
rect 978 1198 1012 1232
rect 1046 1198 1080 1232
rect 1114 1198 1148 1232
rect 1182 1198 1216 1232
rect 1250 1198 1284 1232
rect 1318 1198 1352 1232
rect 1386 1198 1420 1232
rect 1454 1198 1488 1232
rect 570 1042 604 1076
rect 638 1042 672 1076
rect 706 1042 740 1076
rect 774 1042 808 1076
rect 842 1042 876 1076
rect 910 1042 944 1076
rect 978 1042 1012 1076
rect 1046 1042 1080 1076
rect 1114 1042 1148 1076
rect 1182 1042 1216 1076
rect 1250 1042 1284 1076
rect 1318 1042 1352 1076
rect 1386 1042 1420 1076
rect 1454 1042 1488 1076
rect 570 886 604 920
rect 638 886 672 920
rect 706 886 740 920
rect 774 886 808 920
rect 842 886 876 920
rect 910 886 944 920
rect 978 886 1012 920
rect 1046 886 1080 920
rect 1114 886 1148 920
rect 1182 886 1216 920
rect 1250 886 1284 920
rect 1318 886 1352 920
rect 1386 886 1420 920
rect 1454 886 1488 920
rect 570 756 604 790
rect 638 756 672 790
rect 706 756 740 790
rect 774 756 808 790
rect 842 756 876 790
rect 910 756 944 790
rect 978 756 1012 790
rect 1046 756 1080 790
rect 1114 756 1148 790
rect 1182 756 1216 790
rect 1250 756 1284 790
rect 1318 756 1352 790
rect 1386 756 1420 790
rect 1454 756 1488 790
rect 570 600 604 634
rect 638 600 672 634
rect 706 600 740 634
rect 774 600 808 634
rect 842 600 876 634
rect 910 600 944 634
rect 978 600 1012 634
rect 1046 600 1080 634
rect 1114 600 1148 634
rect 1182 600 1216 634
rect 1250 600 1284 634
rect 1318 600 1352 634
rect 1386 600 1420 634
rect 1454 600 1488 634
rect 570 444 604 478
rect 638 444 672 478
rect 706 444 740 478
rect 774 444 808 478
rect 842 444 876 478
rect 910 444 944 478
rect 978 444 1012 478
rect 1046 444 1080 478
rect 1114 444 1148 478
rect 1182 444 1216 478
rect 1250 444 1284 478
rect 1318 444 1352 478
rect 1386 444 1420 478
rect 1454 444 1488 478
rect 2405 1224 2439 1258
rect 2473 1224 2507 1258
rect 2541 1224 2575 1258
rect 2609 1224 2643 1258
rect 2677 1224 2711 1258
rect 2745 1224 2779 1258
rect 2813 1224 2847 1258
rect 2881 1224 2915 1258
rect 2949 1224 2983 1258
rect 3017 1224 3051 1258
rect 3085 1224 3119 1258
rect 3153 1224 3187 1258
rect 3221 1224 3255 1258
rect 3289 1224 3323 1258
rect 3357 1224 3391 1258
rect 3425 1224 3459 1258
rect 3493 1224 3527 1258
rect 3561 1224 3595 1258
rect 3629 1224 3663 1258
rect 3697 1224 3731 1258
rect 3765 1224 3799 1258
rect 3833 1224 3867 1258
rect 3901 1224 3935 1258
rect 3969 1224 4003 1258
rect 4037 1224 4071 1258
rect 4105 1224 4139 1258
rect 4173 1224 4207 1258
rect 4241 1224 4275 1258
rect 4309 1224 4343 1258
rect 4549 1224 4583 1258
rect 4617 1224 4651 1258
rect 4685 1224 4719 1258
rect 4753 1224 4787 1258
rect 4821 1224 4855 1258
rect 4889 1224 4923 1258
rect 4957 1224 4991 1258
rect 5025 1224 5059 1258
rect 5093 1224 5127 1258
rect 5161 1224 5195 1258
rect 5229 1224 5263 1258
rect 5297 1224 5331 1258
rect 5365 1224 5399 1258
rect 5433 1224 5467 1258
rect 5501 1224 5535 1258
rect 5569 1224 5603 1258
rect 5637 1224 5671 1258
rect 5705 1224 5739 1258
rect 5773 1224 5807 1258
rect 5841 1224 5875 1258
rect 5909 1224 5943 1258
rect 5977 1224 6011 1258
rect 6045 1224 6079 1258
rect 6113 1224 6147 1258
rect 6181 1224 6215 1258
rect 6249 1224 6283 1258
rect 6317 1224 6351 1258
rect 6385 1224 6419 1258
rect 6453 1224 6487 1258
rect 2405 1068 2439 1102
rect 2473 1068 2507 1102
rect 2541 1068 2575 1102
rect 2609 1068 2643 1102
rect 2677 1068 2711 1102
rect 2745 1068 2779 1102
rect 2813 1068 2847 1102
rect 2881 1068 2915 1102
rect 2949 1068 2983 1102
rect 3017 1068 3051 1102
rect 3085 1068 3119 1102
rect 3153 1068 3187 1102
rect 3221 1068 3255 1102
rect 3289 1068 3323 1102
rect 3357 1068 3391 1102
rect 3425 1068 3459 1102
rect 3493 1068 3527 1102
rect 3561 1068 3595 1102
rect 3629 1068 3663 1102
rect 3697 1068 3731 1102
rect 3765 1068 3799 1102
rect 3833 1068 3867 1102
rect 3901 1068 3935 1102
rect 3969 1068 4003 1102
rect 4037 1068 4071 1102
rect 4105 1068 4139 1102
rect 4173 1068 4207 1102
rect 4241 1068 4275 1102
rect 4309 1068 4343 1102
rect 4549 1068 4583 1102
rect 4617 1068 4651 1102
rect 4685 1068 4719 1102
rect 4753 1068 4787 1102
rect 4821 1068 4855 1102
rect 4889 1068 4923 1102
rect 4957 1068 4991 1102
rect 5025 1068 5059 1102
rect 5093 1068 5127 1102
rect 5161 1068 5195 1102
rect 5229 1068 5263 1102
rect 5297 1068 5331 1102
rect 5365 1068 5399 1102
rect 5433 1068 5467 1102
rect 5501 1068 5535 1102
rect 5569 1068 5603 1102
rect 5637 1068 5671 1102
rect 5705 1068 5739 1102
rect 5773 1068 5807 1102
rect 5841 1068 5875 1102
rect 5909 1068 5943 1102
rect 5977 1068 6011 1102
rect 6045 1068 6079 1102
rect 6113 1068 6147 1102
rect 6181 1068 6215 1102
rect 6249 1068 6283 1102
rect 6317 1068 6351 1102
rect 6385 1068 6419 1102
rect 6453 1068 6487 1102
rect 2405 912 2439 946
rect 2473 912 2507 946
rect 2541 912 2575 946
rect 2609 912 2643 946
rect 2677 912 2711 946
rect 2745 912 2779 946
rect 2813 912 2847 946
rect 2881 912 2915 946
rect 2949 912 2983 946
rect 3017 912 3051 946
rect 3085 912 3119 946
rect 3153 912 3187 946
rect 3221 912 3255 946
rect 3289 912 3323 946
rect 3357 912 3391 946
rect 3425 912 3459 946
rect 3493 912 3527 946
rect 3561 912 3595 946
rect 3629 912 3663 946
rect 3697 912 3731 946
rect 3765 912 3799 946
rect 3833 912 3867 946
rect 3901 912 3935 946
rect 3969 912 4003 946
rect 4037 912 4071 946
rect 4105 912 4139 946
rect 4173 912 4207 946
rect 4241 912 4275 946
rect 4309 912 4343 946
rect 4549 912 4583 946
rect 4617 912 4651 946
rect 4685 912 4719 946
rect 4753 912 4787 946
rect 4821 912 4855 946
rect 4889 912 4923 946
rect 4957 912 4991 946
rect 5025 912 5059 946
rect 5093 912 5127 946
rect 5161 912 5195 946
rect 5229 912 5263 946
rect 5297 912 5331 946
rect 5365 912 5399 946
rect 5433 912 5467 946
rect 5501 912 5535 946
rect 5569 912 5603 946
rect 5637 912 5671 946
rect 5705 912 5739 946
rect 5773 912 5807 946
rect 5841 912 5875 946
rect 5909 912 5943 946
rect 5977 912 6011 946
rect 6045 912 6079 946
rect 6113 912 6147 946
rect 6181 912 6215 946
rect 6249 912 6283 946
rect 6317 912 6351 946
rect 6385 912 6419 946
rect 6453 912 6487 946
rect 2405 756 2439 790
rect 2473 756 2507 790
rect 2541 756 2575 790
rect 2609 756 2643 790
rect 2677 756 2711 790
rect 2745 756 2779 790
rect 2813 756 2847 790
rect 2881 756 2915 790
rect 2949 756 2983 790
rect 3017 756 3051 790
rect 3085 756 3119 790
rect 3153 756 3187 790
rect 3221 756 3255 790
rect 3289 756 3323 790
rect 3357 756 3391 790
rect 3425 756 3459 790
rect 3493 756 3527 790
rect 3561 756 3595 790
rect 3629 756 3663 790
rect 3697 756 3731 790
rect 3765 756 3799 790
rect 3833 756 3867 790
rect 3901 756 3935 790
rect 3969 756 4003 790
rect 4037 756 4071 790
rect 4105 756 4139 790
rect 4173 756 4207 790
rect 4241 756 4275 790
rect 4309 756 4343 790
rect 4549 756 4583 790
rect 4617 756 4651 790
rect 4685 756 4719 790
rect 4753 756 4787 790
rect 4821 756 4855 790
rect 4889 756 4923 790
rect 4957 756 4991 790
rect 5025 756 5059 790
rect 5093 756 5127 790
rect 5161 756 5195 790
rect 5229 756 5263 790
rect 5297 756 5331 790
rect 5365 756 5399 790
rect 5433 756 5467 790
rect 5501 756 5535 790
rect 5569 756 5603 790
rect 5637 756 5671 790
rect 5705 756 5739 790
rect 5773 756 5807 790
rect 5841 756 5875 790
rect 5909 756 5943 790
rect 5977 756 6011 790
rect 6045 756 6079 790
rect 6113 756 6147 790
rect 6181 756 6215 790
rect 6249 756 6283 790
rect 6317 756 6351 790
rect 6385 756 6419 790
rect 6453 756 6487 790
rect 2405 600 2439 634
rect 2473 600 2507 634
rect 2541 600 2575 634
rect 2609 600 2643 634
rect 2677 600 2711 634
rect 2745 600 2779 634
rect 2813 600 2847 634
rect 2881 600 2915 634
rect 2949 600 2983 634
rect 3017 600 3051 634
rect 3085 600 3119 634
rect 3153 600 3187 634
rect 3221 600 3255 634
rect 3289 600 3323 634
rect 3357 600 3391 634
rect 3425 600 3459 634
rect 3493 600 3527 634
rect 3561 600 3595 634
rect 3629 600 3663 634
rect 3697 600 3731 634
rect 3765 600 3799 634
rect 3833 600 3867 634
rect 3901 600 3935 634
rect 3969 600 4003 634
rect 4037 600 4071 634
rect 4105 600 4139 634
rect 4173 600 4207 634
rect 4241 600 4275 634
rect 4309 600 4343 634
rect 4549 600 4583 634
rect 4617 600 4651 634
rect 4685 600 4719 634
rect 4753 600 4787 634
rect 4821 600 4855 634
rect 4889 600 4923 634
rect 4957 600 4991 634
rect 5025 600 5059 634
rect 5093 600 5127 634
rect 5161 600 5195 634
rect 5229 600 5263 634
rect 5297 600 5331 634
rect 5365 600 5399 634
rect 5433 600 5467 634
rect 5501 600 5535 634
rect 5569 600 5603 634
rect 5637 600 5671 634
rect 5705 600 5739 634
rect 5773 600 5807 634
rect 5841 600 5875 634
rect 5909 600 5943 634
rect 5977 600 6011 634
rect 6045 600 6079 634
rect 6113 600 6147 634
rect 6181 600 6215 634
rect 6249 600 6283 634
rect 6317 600 6351 634
rect 6385 600 6419 634
rect 6453 600 6487 634
rect 2405 444 2439 478
rect 2473 444 2507 478
rect 2541 444 2575 478
rect 2609 444 2643 478
rect 2677 444 2711 478
rect 2745 444 2779 478
rect 2813 444 2847 478
rect 2881 444 2915 478
rect 2949 444 2983 478
rect 3017 444 3051 478
rect 3085 444 3119 478
rect 3153 444 3187 478
rect 3221 444 3255 478
rect 3289 444 3323 478
rect 3357 444 3391 478
rect 3425 444 3459 478
rect 3493 444 3527 478
rect 3561 444 3595 478
rect 3629 444 3663 478
rect 3697 444 3731 478
rect 3765 444 3799 478
rect 3833 444 3867 478
rect 3901 444 3935 478
rect 3969 444 4003 478
rect 4037 444 4071 478
rect 4105 444 4139 478
rect 4173 444 4207 478
rect 4241 444 4275 478
rect 4309 444 4343 478
rect 4549 444 4583 478
rect 4617 444 4651 478
rect 4685 444 4719 478
rect 4753 444 4787 478
rect 4821 444 4855 478
rect 4889 444 4923 478
rect 4957 444 4991 478
rect 5025 444 5059 478
rect 5093 444 5127 478
rect 5161 444 5195 478
rect 5229 444 5263 478
rect 5297 444 5331 478
rect 5365 444 5399 478
rect 5433 444 5467 478
rect 5501 444 5535 478
rect 5569 444 5603 478
rect 5637 444 5671 478
rect 5705 444 5739 478
rect 5773 444 5807 478
rect 5841 444 5875 478
rect 5909 444 5943 478
rect 5977 444 6011 478
rect 6045 444 6079 478
rect 6113 444 6147 478
rect 6181 444 6215 478
rect 6249 444 6283 478
rect 6317 444 6351 478
rect 6385 444 6419 478
rect 6453 444 6487 478
rect 7462 1224 7496 1258
rect 7530 1224 7564 1258
rect 7598 1224 7632 1258
rect 7666 1224 7700 1258
rect 7734 1224 7768 1258
rect 7802 1224 7836 1258
rect 7870 1224 7904 1258
rect 7938 1224 7972 1258
rect 8006 1224 8040 1258
rect 8074 1224 8108 1258
rect 8142 1224 8176 1258
rect 8210 1224 8244 1258
rect 8278 1224 8312 1258
rect 8346 1224 8380 1258
rect 8414 1224 8448 1258
rect 8482 1224 8516 1258
rect 8550 1224 8584 1258
rect 8618 1224 8652 1258
rect 8686 1224 8720 1258
rect 8754 1224 8788 1258
rect 8822 1224 8856 1258
rect 8890 1224 8924 1258
rect 8958 1224 8992 1258
rect 9026 1224 9060 1258
rect 9094 1224 9128 1258
rect 9162 1224 9196 1258
rect 9230 1224 9264 1258
rect 9298 1224 9332 1258
rect 9366 1224 9400 1258
rect 9568 1224 9602 1258
rect 9636 1224 9670 1258
rect 9704 1224 9738 1258
rect 9772 1224 9806 1258
rect 9840 1224 9874 1258
rect 9908 1224 9942 1258
rect 9976 1224 10010 1258
rect 10044 1224 10078 1258
rect 10112 1224 10146 1258
rect 10180 1224 10214 1258
rect 10248 1224 10282 1258
rect 10316 1224 10350 1258
rect 10384 1224 10418 1258
rect 10452 1224 10486 1258
rect 10520 1224 10554 1258
rect 10588 1224 10622 1258
rect 10656 1224 10690 1258
rect 10724 1224 10758 1258
rect 10792 1224 10826 1258
rect 10860 1224 10894 1258
rect 10928 1224 10962 1258
rect 10996 1224 11030 1258
rect 11064 1224 11098 1258
rect 11132 1224 11166 1258
rect 11200 1224 11234 1258
rect 11268 1224 11302 1258
rect 11336 1224 11370 1258
rect 11404 1224 11438 1258
rect 11472 1224 11506 1258
rect 7462 1068 7496 1102
rect 7530 1068 7564 1102
rect 7598 1068 7632 1102
rect 7666 1068 7700 1102
rect 7734 1068 7768 1102
rect 7802 1068 7836 1102
rect 7870 1068 7904 1102
rect 7938 1068 7972 1102
rect 8006 1068 8040 1102
rect 8074 1068 8108 1102
rect 8142 1068 8176 1102
rect 8210 1068 8244 1102
rect 8278 1068 8312 1102
rect 8346 1068 8380 1102
rect 8414 1068 8448 1102
rect 8482 1068 8516 1102
rect 8550 1068 8584 1102
rect 8618 1068 8652 1102
rect 8686 1068 8720 1102
rect 8754 1068 8788 1102
rect 8822 1068 8856 1102
rect 8890 1068 8924 1102
rect 8958 1068 8992 1102
rect 9026 1068 9060 1102
rect 9094 1068 9128 1102
rect 9162 1068 9196 1102
rect 9230 1068 9264 1102
rect 9298 1068 9332 1102
rect 9366 1068 9400 1102
rect 9568 1068 9602 1102
rect 9636 1068 9670 1102
rect 9704 1068 9738 1102
rect 9772 1068 9806 1102
rect 9840 1068 9874 1102
rect 9908 1068 9942 1102
rect 9976 1068 10010 1102
rect 10044 1068 10078 1102
rect 10112 1068 10146 1102
rect 10180 1068 10214 1102
rect 10248 1068 10282 1102
rect 10316 1068 10350 1102
rect 10384 1068 10418 1102
rect 10452 1068 10486 1102
rect 10520 1068 10554 1102
rect 10588 1068 10622 1102
rect 10656 1068 10690 1102
rect 10724 1068 10758 1102
rect 10792 1068 10826 1102
rect 10860 1068 10894 1102
rect 10928 1068 10962 1102
rect 10996 1068 11030 1102
rect 11064 1068 11098 1102
rect 11132 1068 11166 1102
rect 11200 1068 11234 1102
rect 11268 1068 11302 1102
rect 11336 1068 11370 1102
rect 11404 1068 11438 1102
rect 11472 1068 11506 1102
rect 7462 912 7496 946
rect 7530 912 7564 946
rect 7598 912 7632 946
rect 7666 912 7700 946
rect 7734 912 7768 946
rect 7802 912 7836 946
rect 7870 912 7904 946
rect 7938 912 7972 946
rect 8006 912 8040 946
rect 8074 912 8108 946
rect 8142 912 8176 946
rect 8210 912 8244 946
rect 8278 912 8312 946
rect 8346 912 8380 946
rect 8414 912 8448 946
rect 8482 912 8516 946
rect 8550 912 8584 946
rect 8618 912 8652 946
rect 8686 912 8720 946
rect 8754 912 8788 946
rect 8822 912 8856 946
rect 8890 912 8924 946
rect 8958 912 8992 946
rect 9026 912 9060 946
rect 9094 912 9128 946
rect 9162 912 9196 946
rect 9230 912 9264 946
rect 9298 912 9332 946
rect 9366 912 9400 946
rect 9568 912 9602 946
rect 9636 912 9670 946
rect 9704 912 9738 946
rect 9772 912 9806 946
rect 9840 912 9874 946
rect 9908 912 9942 946
rect 9976 912 10010 946
rect 10044 912 10078 946
rect 10112 912 10146 946
rect 10180 912 10214 946
rect 10248 912 10282 946
rect 10316 912 10350 946
rect 10384 912 10418 946
rect 10452 912 10486 946
rect 10520 912 10554 946
rect 10588 912 10622 946
rect 10656 912 10690 946
rect 10724 912 10758 946
rect 10792 912 10826 946
rect 10860 912 10894 946
rect 10928 912 10962 946
rect 10996 912 11030 946
rect 11064 912 11098 946
rect 11132 912 11166 946
rect 11200 912 11234 946
rect 11268 912 11302 946
rect 11336 912 11370 946
rect 11404 912 11438 946
rect 11472 912 11506 946
rect 7462 756 7496 790
rect 7530 756 7564 790
rect 7598 756 7632 790
rect 7666 756 7700 790
rect 7734 756 7768 790
rect 7802 756 7836 790
rect 7870 756 7904 790
rect 7938 756 7972 790
rect 8006 756 8040 790
rect 8074 756 8108 790
rect 8142 756 8176 790
rect 8210 756 8244 790
rect 8278 756 8312 790
rect 8346 756 8380 790
rect 8414 756 8448 790
rect 8482 756 8516 790
rect 8550 756 8584 790
rect 8618 756 8652 790
rect 8686 756 8720 790
rect 8754 756 8788 790
rect 8822 756 8856 790
rect 8890 756 8924 790
rect 8958 756 8992 790
rect 9026 756 9060 790
rect 9094 756 9128 790
rect 9162 756 9196 790
rect 9230 756 9264 790
rect 9298 756 9332 790
rect 9366 756 9400 790
rect 9568 756 9602 790
rect 9636 756 9670 790
rect 9704 756 9738 790
rect 9772 756 9806 790
rect 9840 756 9874 790
rect 9908 756 9942 790
rect 9976 756 10010 790
rect 10044 756 10078 790
rect 10112 756 10146 790
rect 10180 756 10214 790
rect 10248 756 10282 790
rect 10316 756 10350 790
rect 10384 756 10418 790
rect 10452 756 10486 790
rect 10520 756 10554 790
rect 10588 756 10622 790
rect 10656 756 10690 790
rect 10724 756 10758 790
rect 10792 756 10826 790
rect 10860 756 10894 790
rect 10928 756 10962 790
rect 10996 756 11030 790
rect 11064 756 11098 790
rect 11132 756 11166 790
rect 11200 756 11234 790
rect 11268 756 11302 790
rect 11336 756 11370 790
rect 11404 756 11438 790
rect 11472 756 11506 790
rect 7462 600 7496 634
rect 7530 600 7564 634
rect 7598 600 7632 634
rect 7666 600 7700 634
rect 7734 600 7768 634
rect 7802 600 7836 634
rect 7870 600 7904 634
rect 7938 600 7972 634
rect 8006 600 8040 634
rect 8074 600 8108 634
rect 8142 600 8176 634
rect 8210 600 8244 634
rect 8278 600 8312 634
rect 8346 600 8380 634
rect 8414 600 8448 634
rect 8482 600 8516 634
rect 8550 600 8584 634
rect 8618 600 8652 634
rect 8686 600 8720 634
rect 8754 600 8788 634
rect 8822 600 8856 634
rect 8890 600 8924 634
rect 8958 600 8992 634
rect 9026 600 9060 634
rect 9094 600 9128 634
rect 9162 600 9196 634
rect 9230 600 9264 634
rect 9298 600 9332 634
rect 9366 600 9400 634
rect 9568 600 9602 634
rect 9636 600 9670 634
rect 9704 600 9738 634
rect 9772 600 9806 634
rect 9840 600 9874 634
rect 9908 600 9942 634
rect 9976 600 10010 634
rect 10044 600 10078 634
rect 10112 600 10146 634
rect 10180 600 10214 634
rect 10248 600 10282 634
rect 10316 600 10350 634
rect 10384 600 10418 634
rect 10452 600 10486 634
rect 10520 600 10554 634
rect 10588 600 10622 634
rect 10656 600 10690 634
rect 10724 600 10758 634
rect 10792 600 10826 634
rect 10860 600 10894 634
rect 10928 600 10962 634
rect 10996 600 11030 634
rect 11064 600 11098 634
rect 11132 600 11166 634
rect 11200 600 11234 634
rect 11268 600 11302 634
rect 11336 600 11370 634
rect 11404 600 11438 634
rect 11472 600 11506 634
rect 7462 444 7496 478
rect 7530 444 7564 478
rect 7598 444 7632 478
rect 7666 444 7700 478
rect 7734 444 7768 478
rect 7802 444 7836 478
rect 7870 444 7904 478
rect 7938 444 7972 478
rect 8006 444 8040 478
rect 8074 444 8108 478
rect 8142 444 8176 478
rect 8210 444 8244 478
rect 8278 444 8312 478
rect 8346 444 8380 478
rect 8414 444 8448 478
rect 8482 444 8516 478
rect 8550 444 8584 478
rect 8618 444 8652 478
rect 8686 444 8720 478
rect 8754 444 8788 478
rect 8822 444 8856 478
rect 8890 444 8924 478
rect 8958 444 8992 478
rect 9026 444 9060 478
rect 9094 444 9128 478
rect 9162 444 9196 478
rect 9230 444 9264 478
rect 9298 444 9332 478
rect 9366 444 9400 478
rect 9568 444 9602 478
rect 9636 444 9670 478
rect 9704 444 9738 478
rect 9772 444 9806 478
rect 9840 444 9874 478
rect 9908 444 9942 478
rect 9976 444 10010 478
rect 10044 444 10078 478
rect 10112 444 10146 478
rect 10180 444 10214 478
rect 10248 444 10282 478
rect 10316 444 10350 478
rect 10384 444 10418 478
rect 10452 444 10486 478
rect 10520 444 10554 478
rect 10588 444 10622 478
rect 10656 444 10690 478
rect 10724 444 10758 478
rect 10792 444 10826 478
rect 10860 444 10894 478
rect 10928 444 10962 478
rect 10996 444 11030 478
rect 11064 444 11098 478
rect 11132 444 11166 478
rect 11200 444 11234 478
rect 11268 444 11302 478
rect 11336 444 11370 478
rect 11404 444 11438 478
rect 11472 444 11506 478
<< mvpdiffc >>
rect 5866 -1304 5900 -1270
rect 5934 -1304 5968 -1270
rect 6002 -1304 6036 -1270
rect 6070 -1304 6104 -1270
rect 6138 -1304 6172 -1270
rect 6206 -1304 6240 -1270
rect 6274 -1304 6308 -1270
rect 6342 -1304 6376 -1270
rect 6410 -1304 6444 -1270
rect 6478 -1304 6512 -1270
rect 6546 -1304 6580 -1270
rect 6614 -1304 6648 -1270
rect 6682 -1304 6716 -1270
rect 6750 -1304 6784 -1270
rect 6818 -1304 6852 -1270
rect 6886 -1304 6920 -1270
rect 6954 -1304 6988 -1270
rect 7022 -1304 7056 -1270
rect 7090 -1304 7124 -1270
rect 7158 -1304 7192 -1270
rect 7226 -1304 7260 -1270
rect 7294 -1304 7328 -1270
rect 7362 -1304 7396 -1270
rect 7430 -1304 7464 -1270
rect 7498 -1304 7532 -1270
rect 7566 -1304 7600 -1270
rect 7634 -1304 7668 -1270
rect 7702 -1304 7736 -1270
rect 7770 -1304 7804 -1270
rect 5866 -1460 5900 -1426
rect 5934 -1460 5968 -1426
rect 6002 -1460 6036 -1426
rect 6070 -1460 6104 -1426
rect 6138 -1460 6172 -1426
rect 6206 -1460 6240 -1426
rect 6274 -1460 6308 -1426
rect 6342 -1460 6376 -1426
rect 6410 -1460 6444 -1426
rect 6478 -1460 6512 -1426
rect 6546 -1460 6580 -1426
rect 6614 -1460 6648 -1426
rect 6682 -1460 6716 -1426
rect 6750 -1460 6784 -1426
rect 6818 -1460 6852 -1426
rect 6886 -1460 6920 -1426
rect 6954 -1460 6988 -1426
rect 7022 -1460 7056 -1426
rect 7090 -1460 7124 -1426
rect 7158 -1460 7192 -1426
rect 7226 -1460 7260 -1426
rect 7294 -1460 7328 -1426
rect 7362 -1460 7396 -1426
rect 7430 -1460 7464 -1426
rect 7498 -1460 7532 -1426
rect 7566 -1460 7600 -1426
rect 7634 -1460 7668 -1426
rect 7702 -1460 7736 -1426
rect 7770 -1460 7804 -1426
rect 5866 -1616 5900 -1582
rect 5934 -1616 5968 -1582
rect 6002 -1616 6036 -1582
rect 6070 -1616 6104 -1582
rect 6138 -1616 6172 -1582
rect 6206 -1616 6240 -1582
rect 6274 -1616 6308 -1582
rect 6342 -1616 6376 -1582
rect 6410 -1616 6444 -1582
rect 6478 -1616 6512 -1582
rect 6546 -1616 6580 -1582
rect 6614 -1616 6648 -1582
rect 6682 -1616 6716 -1582
rect 6750 -1616 6784 -1582
rect 6818 -1616 6852 -1582
rect 6886 -1616 6920 -1582
rect 6954 -1616 6988 -1582
rect 7022 -1616 7056 -1582
rect 7090 -1616 7124 -1582
rect 7158 -1616 7192 -1582
rect 7226 -1616 7260 -1582
rect 7294 -1616 7328 -1582
rect 7362 -1616 7396 -1582
rect 7430 -1616 7464 -1582
rect 7498 -1616 7532 -1582
rect 7566 -1616 7600 -1582
rect 7634 -1616 7668 -1582
rect 7702 -1616 7736 -1582
rect 7770 -1616 7804 -1582
rect 5866 -1772 5900 -1738
rect 5934 -1772 5968 -1738
rect 6002 -1772 6036 -1738
rect 6070 -1772 6104 -1738
rect 6138 -1772 6172 -1738
rect 6206 -1772 6240 -1738
rect 6274 -1772 6308 -1738
rect 6342 -1772 6376 -1738
rect 6410 -1772 6444 -1738
rect 6478 -1772 6512 -1738
rect 6546 -1772 6580 -1738
rect 6614 -1772 6648 -1738
rect 6682 -1772 6716 -1738
rect 6750 -1772 6784 -1738
rect 6818 -1772 6852 -1738
rect 6886 -1772 6920 -1738
rect 6954 -1772 6988 -1738
rect 7022 -1772 7056 -1738
rect 7090 -1772 7124 -1738
rect 7158 -1772 7192 -1738
rect 7226 -1772 7260 -1738
rect 7294 -1772 7328 -1738
rect 7362 -1772 7396 -1738
rect 7430 -1772 7464 -1738
rect 7498 -1772 7532 -1738
rect 7566 -1772 7600 -1738
rect 7634 -1772 7668 -1738
rect 7702 -1772 7736 -1738
rect 7770 -1772 7804 -1738
rect 5866 -1928 5900 -1894
rect 5934 -1928 5968 -1894
rect 6002 -1928 6036 -1894
rect 6070 -1928 6104 -1894
rect 6138 -1928 6172 -1894
rect 6206 -1928 6240 -1894
rect 6274 -1928 6308 -1894
rect 6342 -1928 6376 -1894
rect 6410 -1928 6444 -1894
rect 6478 -1928 6512 -1894
rect 6546 -1928 6580 -1894
rect 6614 -1928 6648 -1894
rect 6682 -1928 6716 -1894
rect 6750 -1928 6784 -1894
rect 6818 -1928 6852 -1894
rect 6886 -1928 6920 -1894
rect 6954 -1928 6988 -1894
rect 7022 -1928 7056 -1894
rect 7090 -1928 7124 -1894
rect 7158 -1928 7192 -1894
rect 7226 -1928 7260 -1894
rect 7294 -1928 7328 -1894
rect 7362 -1928 7396 -1894
rect 7430 -1928 7464 -1894
rect 7498 -1928 7532 -1894
rect 7566 -1928 7600 -1894
rect 7634 -1928 7668 -1894
rect 7702 -1928 7736 -1894
rect 7770 -1928 7804 -1894
<< mvpsubdiff >>
rect 357 1351 1709 1354
rect 357 1317 458 1351
rect 492 1317 526 1351
rect 560 1317 594 1351
rect 628 1317 662 1351
rect 696 1317 730 1351
rect 764 1317 798 1351
rect 832 1317 866 1351
rect 900 1317 934 1351
rect 968 1317 1002 1351
rect 1036 1317 1131 1351
rect 1165 1317 1199 1351
rect 1233 1317 1267 1351
rect 1301 1317 1335 1351
rect 1369 1317 1403 1351
rect 1437 1317 1471 1351
rect 1505 1317 1539 1351
rect 1573 1317 1607 1351
rect 1641 1317 1709 1351
rect 357 1314 1709 1317
rect 357 1286 397 1314
rect 357 1252 360 1286
rect 394 1252 397 1286
rect 357 1218 397 1252
rect 357 1184 360 1218
rect 394 1184 397 1218
rect 357 1150 397 1184
rect 357 1116 360 1150
rect 394 1116 397 1150
rect 357 1082 397 1116
rect 357 1048 360 1082
rect 394 1048 397 1082
rect 357 1014 397 1048
rect 357 980 360 1014
rect 394 980 397 1014
rect 357 946 397 980
rect 357 912 360 946
rect 394 912 397 946
rect 357 878 397 912
rect 357 844 360 878
rect 394 844 397 878
rect 357 810 397 844
rect 357 776 360 810
rect 394 776 397 810
rect 357 742 397 776
rect 357 708 360 742
rect 394 708 397 742
rect 357 674 397 708
rect 357 640 360 674
rect 394 640 397 674
rect 357 606 397 640
rect 357 572 360 606
rect 394 572 397 606
rect 357 538 397 572
rect 1669 1240 1709 1314
rect 1669 1206 1672 1240
rect 1706 1206 1709 1240
rect 1669 1172 1709 1206
rect 1669 1138 1672 1172
rect 1706 1138 1709 1172
rect 1669 1104 1709 1138
rect 1669 1070 1672 1104
rect 1706 1070 1709 1104
rect 1669 1036 1709 1070
rect 1669 1002 1672 1036
rect 1706 1002 1709 1036
rect 1669 968 1709 1002
rect 1669 934 1672 968
rect 1706 934 1709 968
rect 1669 900 1709 934
rect 1669 866 1672 900
rect 1706 866 1709 900
rect 1669 832 1709 866
rect 1669 798 1672 832
rect 1706 798 1709 832
rect 1669 764 1709 798
rect 1669 730 1672 764
rect 1706 730 1709 764
rect 1669 696 1709 730
rect 1669 662 1672 696
rect 1706 662 1709 696
rect 1669 628 1709 662
rect 1669 594 1672 628
rect 1706 594 1709 628
rect 357 504 360 538
rect 394 504 397 538
rect 357 470 397 504
rect 1669 560 1709 594
rect 1669 526 1672 560
rect 1706 526 1709 560
rect 1669 492 1709 526
rect 357 436 360 470
rect 394 436 397 470
rect 1669 458 1672 492
rect 1706 458 1709 492
rect 357 362 397 436
rect 1669 424 1709 458
rect 1669 390 1672 424
rect 1706 390 1709 424
rect 1669 362 1709 390
rect 357 359 1709 362
rect 357 325 425 359
rect 459 325 493 359
rect 527 325 561 359
rect 595 325 629 359
rect 663 325 697 359
rect 731 325 765 359
rect 799 325 833 359
rect 867 325 901 359
rect 935 325 969 359
rect 1003 325 1037 359
rect 1071 325 1105 359
rect 1139 325 1173 359
rect 1207 325 1241 359
rect 1275 325 1309 359
rect 1343 325 1377 359
rect 1411 325 1445 359
rect 1479 325 1513 359
rect 1547 325 1581 359
rect 1615 325 1709 359
rect 357 322 1709 325
rect 2192 1377 6700 1380
rect 2192 1343 2287 1377
rect 2321 1343 2355 1377
rect 2389 1343 2423 1377
rect 2457 1343 2491 1377
rect 2525 1343 2559 1377
rect 2593 1343 2627 1377
rect 2661 1343 2695 1377
rect 2729 1343 2763 1377
rect 2797 1343 2831 1377
rect 2865 1343 2899 1377
rect 2933 1343 2967 1377
rect 3001 1343 3035 1377
rect 3069 1343 3103 1377
rect 3137 1343 3171 1377
rect 3205 1343 3239 1377
rect 3273 1343 3307 1377
rect 3341 1343 3375 1377
rect 3409 1343 3443 1377
rect 3477 1343 3511 1377
rect 3545 1343 3579 1377
rect 3613 1343 3647 1377
rect 3681 1343 3715 1377
rect 3749 1343 3783 1377
rect 3817 1343 3851 1377
rect 3885 1343 3919 1377
rect 3953 1343 3987 1377
rect 4021 1343 4055 1377
rect 4089 1343 4123 1377
rect 4157 1343 4191 1377
rect 4225 1343 4259 1377
rect 4293 1343 4327 1377
rect 4361 1343 4395 1377
rect 4429 1343 4558 1377
rect 4592 1343 4626 1377
rect 4660 1343 4694 1377
rect 4728 1343 4762 1377
rect 4796 1343 4830 1377
rect 4864 1343 4898 1377
rect 4932 1343 4966 1377
rect 5000 1343 5034 1377
rect 5068 1343 5102 1377
rect 5136 1343 5170 1377
rect 5204 1343 5238 1377
rect 5272 1343 5306 1377
rect 5340 1343 5374 1377
rect 5408 1343 5442 1377
rect 5476 1343 5510 1377
rect 5544 1343 5578 1377
rect 5612 1343 5646 1377
rect 5680 1343 5714 1377
rect 5748 1343 5782 1377
rect 5816 1343 5850 1377
rect 5884 1343 5918 1377
rect 5952 1343 5986 1377
rect 6020 1343 6054 1377
rect 6088 1343 6122 1377
rect 6156 1343 6190 1377
rect 6224 1343 6258 1377
rect 6292 1343 6326 1377
rect 6360 1343 6394 1377
rect 6428 1343 6462 1377
rect 6496 1343 6530 1377
rect 6564 1343 6598 1377
rect 6632 1343 6700 1377
rect 2192 1340 6700 1343
rect 2192 1312 2232 1340
rect 2192 1278 2195 1312
rect 2229 1278 2232 1312
rect 2192 1244 2232 1278
rect 6660 1308 6700 1340
rect 6660 1274 6663 1308
rect 6697 1274 6700 1308
rect 2192 1210 2195 1244
rect 2229 1210 2232 1244
rect 6660 1240 6700 1274
rect 2192 1176 2232 1210
rect 2192 1142 2195 1176
rect 2229 1142 2232 1176
rect 2192 1108 2232 1142
rect 2192 1074 2195 1108
rect 2229 1074 2232 1108
rect 2192 1040 2232 1074
rect 2192 1006 2195 1040
rect 2229 1006 2232 1040
rect 2192 972 2232 1006
rect 2192 938 2195 972
rect 2229 938 2232 972
rect 2192 904 2232 938
rect 2192 870 2195 904
rect 2229 870 2232 904
rect 2192 836 2232 870
rect 2192 802 2195 836
rect 2229 802 2232 836
rect 2192 768 2232 802
rect 2192 734 2195 768
rect 2229 734 2232 768
rect 2192 700 2232 734
rect 2192 666 2195 700
rect 2229 666 2232 700
rect 2192 632 2232 666
rect 2192 598 2195 632
rect 2229 598 2232 632
rect 2192 564 2232 598
rect 2192 530 2195 564
rect 2229 530 2232 564
rect 2192 496 2232 530
rect 2192 462 2195 496
rect 2229 462 2232 496
rect 6660 1206 6663 1240
rect 6697 1206 6700 1240
rect 6660 1172 6700 1206
rect 6660 1138 6663 1172
rect 6697 1138 6700 1172
rect 6660 1104 6700 1138
rect 6660 1070 6663 1104
rect 6697 1070 6700 1104
rect 6660 1036 6700 1070
rect 6660 1002 6663 1036
rect 6697 1002 6700 1036
rect 6660 968 6700 1002
rect 6660 934 6663 968
rect 6697 934 6700 968
rect 6660 900 6700 934
rect 6660 866 6663 900
rect 6697 866 6700 900
rect 6660 832 6700 866
rect 6660 798 6663 832
rect 6697 798 6700 832
rect 6660 764 6700 798
rect 6660 730 6663 764
rect 6697 730 6700 764
rect 6660 696 6700 730
rect 6660 662 6663 696
rect 6697 662 6700 696
rect 6660 628 6700 662
rect 6660 594 6663 628
rect 6697 594 6700 628
rect 6660 560 6700 594
rect 6660 526 6663 560
rect 6697 526 6700 560
rect 6660 492 6700 526
rect 2192 428 2232 462
rect 6660 458 6663 492
rect 6697 458 6700 492
rect 2192 394 2195 428
rect 2229 394 2232 428
rect 2192 362 2232 394
rect 6660 424 6700 458
rect 6660 390 6663 424
rect 6697 390 6700 424
rect 6660 362 6700 390
rect 2192 359 6700 362
rect 2192 325 2260 359
rect 2294 325 2328 359
rect 2362 325 2396 359
rect 2430 325 2464 359
rect 2498 325 2532 359
rect 2566 325 2600 359
rect 2634 325 2668 359
rect 2702 325 2736 359
rect 2770 325 2804 359
rect 2838 325 2872 359
rect 2906 325 2940 359
rect 2974 325 3008 359
rect 3042 325 3076 359
rect 3110 325 3144 359
rect 3178 325 3212 359
rect 3246 325 3280 359
rect 3314 325 3348 359
rect 3382 325 3416 359
rect 3450 325 3484 359
rect 3518 325 3552 359
rect 3586 325 3620 359
rect 3654 325 3688 359
rect 3722 325 3756 359
rect 3790 325 3824 359
rect 3858 325 3892 359
rect 3926 325 3960 359
rect 3994 325 4028 359
rect 4062 325 4096 359
rect 4130 325 4164 359
rect 4198 325 4232 359
rect 4266 325 4300 359
rect 4334 325 4368 359
rect 4402 325 4436 359
rect 4470 325 4504 359
rect 4538 325 4572 359
rect 4606 325 4640 359
rect 4674 325 4708 359
rect 4742 325 4776 359
rect 4810 325 4844 359
rect 4878 325 4912 359
rect 4946 325 4980 359
rect 5014 325 5048 359
rect 5082 325 5116 359
rect 5150 325 5184 359
rect 5218 325 5252 359
rect 5286 325 5320 359
rect 5354 325 5388 359
rect 5422 325 5456 359
rect 5490 325 5524 359
rect 5558 325 5592 359
rect 5626 325 5660 359
rect 5694 325 5728 359
rect 5762 325 5796 359
rect 5830 325 5864 359
rect 5898 325 5932 359
rect 5966 325 6000 359
rect 6034 325 6068 359
rect 6102 325 6136 359
rect 6170 325 6204 359
rect 6238 325 6272 359
rect 6306 325 6340 359
rect 6374 325 6408 359
rect 6442 325 6476 359
rect 6510 325 6544 359
rect 6578 325 6700 359
rect 2192 322 6700 325
rect 7196 1377 11718 1380
rect 7196 1343 7264 1377
rect 7298 1343 7332 1377
rect 7366 1343 7400 1377
rect 7434 1343 7468 1377
rect 7502 1343 7536 1377
rect 7570 1343 7604 1377
rect 7638 1343 7672 1377
rect 7706 1343 7740 1377
rect 7774 1343 7808 1377
rect 7842 1343 7876 1377
rect 7910 1343 7944 1377
rect 7978 1343 8012 1377
rect 8046 1343 8080 1377
rect 8114 1343 8148 1377
rect 8182 1343 8216 1377
rect 8250 1343 8284 1377
rect 8318 1343 8352 1377
rect 8386 1343 8420 1377
rect 8454 1343 8488 1377
rect 8522 1343 8556 1377
rect 8590 1343 8624 1377
rect 8658 1343 8692 1377
rect 8726 1343 8760 1377
rect 8794 1343 8828 1377
rect 8862 1343 8896 1377
rect 8930 1343 8964 1377
rect 8998 1343 9032 1377
rect 9066 1343 9100 1377
rect 9134 1343 9168 1377
rect 9202 1343 9236 1377
rect 9270 1343 9304 1377
rect 9338 1343 9372 1377
rect 9406 1343 9500 1377
rect 9534 1343 9568 1377
rect 9602 1343 9636 1377
rect 9670 1343 9704 1377
rect 9738 1343 9772 1377
rect 9806 1343 9840 1377
rect 9874 1343 9908 1377
rect 9942 1343 9976 1377
rect 10010 1343 10044 1377
rect 10078 1343 10112 1377
rect 10146 1343 10180 1377
rect 10214 1343 10248 1377
rect 10282 1343 10316 1377
rect 10350 1343 10384 1377
rect 10418 1343 10452 1377
rect 10486 1343 10520 1377
rect 10554 1343 10588 1377
rect 10622 1343 10656 1377
rect 10690 1343 10724 1377
rect 10758 1343 10792 1377
rect 10826 1343 10860 1377
rect 10894 1343 10928 1377
rect 10962 1343 10996 1377
rect 11030 1343 11064 1377
rect 11098 1343 11132 1377
rect 11166 1343 11200 1377
rect 11234 1343 11268 1377
rect 11302 1343 11336 1377
rect 11370 1343 11404 1377
rect 11438 1343 11472 1377
rect 11506 1343 11540 1377
rect 11574 1343 11608 1377
rect 11642 1343 11718 1377
rect 7196 1340 11718 1343
rect 7196 1308 7236 1340
rect 7196 1274 7199 1308
rect 7233 1274 7236 1308
rect 7196 1240 7236 1274
rect 11678 1312 11718 1340
rect 11678 1278 11681 1312
rect 11715 1278 11718 1312
rect 7196 1206 7199 1240
rect 7233 1206 7236 1240
rect 11678 1244 11718 1278
rect 7196 1172 7236 1206
rect 7196 1138 7199 1172
rect 7233 1138 7236 1172
rect 7196 1104 7236 1138
rect 7196 1070 7199 1104
rect 7233 1070 7236 1104
rect 7196 1036 7236 1070
rect 7196 1002 7199 1036
rect 7233 1002 7236 1036
rect 7196 968 7236 1002
rect 7196 934 7199 968
rect 7233 934 7236 968
rect 7196 900 7236 934
rect 7196 866 7199 900
rect 7233 866 7236 900
rect 7196 832 7236 866
rect 7196 798 7199 832
rect 7233 798 7236 832
rect 7196 764 7236 798
rect 7196 730 7199 764
rect 7233 730 7236 764
rect 7196 696 7236 730
rect 7196 662 7199 696
rect 7233 662 7236 696
rect 7196 628 7236 662
rect 7196 594 7199 628
rect 7233 594 7236 628
rect 7196 560 7236 594
rect 7196 526 7199 560
rect 7233 526 7236 560
rect 7196 492 7236 526
rect 7196 458 7199 492
rect 7233 458 7236 492
rect 11678 1210 11681 1244
rect 11715 1210 11718 1244
rect 11678 1176 11718 1210
rect 11678 1142 11681 1176
rect 11715 1142 11718 1176
rect 11678 1108 11718 1142
rect 11678 1074 11681 1108
rect 11715 1074 11718 1108
rect 11678 1040 11718 1074
rect 11678 1006 11681 1040
rect 11715 1006 11718 1040
rect 11678 972 11718 1006
rect 11678 938 11681 972
rect 11715 938 11718 972
rect 11678 904 11718 938
rect 11678 870 11681 904
rect 11715 870 11718 904
rect 11678 836 11718 870
rect 11678 802 11681 836
rect 11715 802 11718 836
rect 11678 768 11718 802
rect 11678 734 11681 768
rect 11715 734 11718 768
rect 11678 700 11718 734
rect 11678 666 11681 700
rect 11715 666 11718 700
rect 11678 632 11718 666
rect 11678 598 11681 632
rect 11715 598 11718 632
rect 11678 564 11718 598
rect 11678 530 11681 564
rect 11715 530 11718 564
rect 11678 496 11718 530
rect 7196 424 7236 458
rect 11678 462 11681 496
rect 11715 462 11718 496
rect 7196 390 7199 424
rect 7233 390 7236 424
rect 7196 362 7236 390
rect 11678 428 11718 462
rect 11678 394 11681 428
rect 11715 394 11718 428
rect 11678 362 11718 394
rect 7196 359 11718 362
rect 7196 325 7264 359
rect 7298 325 7332 359
rect 7366 325 7400 359
rect 7434 325 7468 359
rect 7502 325 7536 359
rect 7570 325 7604 359
rect 7638 325 7672 359
rect 7706 325 7740 359
rect 7774 325 7808 359
rect 7842 325 7876 359
rect 7910 325 7944 359
rect 7978 325 8012 359
rect 8046 325 8080 359
rect 8114 325 8148 359
rect 8182 325 8216 359
rect 8250 325 8284 359
rect 8318 325 8352 359
rect 8386 325 8420 359
rect 8454 325 8488 359
rect 8522 325 8556 359
rect 8590 325 8624 359
rect 8658 325 8692 359
rect 8726 325 8760 359
rect 8794 325 8828 359
rect 8862 325 8896 359
rect 8930 325 8964 359
rect 8998 325 9032 359
rect 9066 325 9100 359
rect 9134 325 9168 359
rect 9202 325 9236 359
rect 9270 325 9304 359
rect 9338 325 9372 359
rect 9406 325 9440 359
rect 9474 325 9508 359
rect 9542 325 9576 359
rect 9610 325 9644 359
rect 9678 325 9712 359
rect 9746 325 9780 359
rect 9814 325 9848 359
rect 9882 325 9916 359
rect 9950 325 9984 359
rect 10018 325 10052 359
rect 10086 325 10120 359
rect 10154 325 10188 359
rect 10222 325 10256 359
rect 10290 325 10324 359
rect 10358 325 10392 359
rect 10426 325 10460 359
rect 10494 325 10528 359
rect 10562 325 10596 359
rect 10630 325 10664 359
rect 10698 325 10732 359
rect 10766 325 10800 359
rect 10834 325 10868 359
rect 10902 325 10936 359
rect 10970 325 11004 359
rect 11038 325 11072 359
rect 11106 325 11140 359
rect 11174 325 11208 359
rect 11242 325 11276 359
rect 11310 325 11344 359
rect 11378 325 11412 359
rect 11446 325 11480 359
rect 11514 325 11548 359
rect 11582 325 11616 359
rect 11650 325 11718 359
rect 7196 322 11718 325
<< mvnsubdiff >>
rect 63 1534 6986 1636
rect 63 1461 165 1534
rect 1906 1461 2008 1534
rect 165 135 206 169
rect 63 101 206 135
rect 63 67 138 101
rect 172 67 206 101
rect 1872 135 1906 169
rect 6884 1450 6986 1534
rect 6884 169 6986 260
rect 2008 135 2103 169
rect 1872 101 2103 135
rect 1872 67 2035 101
rect 2069 67 2103 101
rect 4653 135 7020 169
rect 7054 135 7089 169
rect 7123 135 7158 169
rect 7192 135 7227 169
rect 7261 135 7296 169
rect 7330 135 7365 169
rect 7399 135 7434 169
rect 7468 135 7503 169
rect 7537 135 7572 169
rect 7606 135 7641 169
rect 7675 135 7710 169
rect 7744 135 7779 169
rect 7813 135 7848 169
rect 7882 135 7917 169
rect 7951 135 7986 169
rect 8020 135 8055 169
rect 8089 135 8124 169
rect 8158 135 8193 169
rect 8227 135 8262 169
rect 8296 135 8331 169
rect 8365 135 8400 169
rect 8434 135 8469 169
rect 8503 135 8538 169
rect 8572 135 8607 169
rect 8641 135 8676 169
rect 8710 135 8745 169
rect 8779 135 8814 169
rect 8848 135 8883 169
rect 8917 135 8952 169
rect 4653 101 8952 135
rect 4653 67 7020 101
rect 7054 67 7089 101
rect 7123 67 7158 101
rect 7192 67 7227 101
rect 7261 67 7296 101
rect 7330 67 7365 101
rect 7399 67 7434 101
rect 7468 67 7503 101
rect 7537 67 7572 101
rect 7606 67 7641 101
rect 7675 67 7710 101
rect 7744 67 7779 101
rect 7813 67 7848 101
rect 7882 67 7917 101
rect 7951 67 7986 101
rect 8020 67 8055 101
rect 8089 67 8124 101
rect 8158 67 8193 101
rect 8227 67 8262 101
rect 8296 67 8331 101
rect 8365 67 8400 101
rect 8434 67 8469 101
rect 8503 67 8538 101
rect 8572 67 8607 101
rect 8641 67 8676 101
rect 8710 67 8745 101
rect 8779 67 8814 101
rect 8848 67 8883 101
rect 8917 67 8952 101
rect 11842 67 11905 169
rect 5617 -1188 5698 -1154
rect 5732 -1188 5766 -1154
rect 5800 -1188 5834 -1154
rect 5868 -1188 5902 -1154
rect 5936 -1188 5970 -1154
rect 6004 -1188 6038 -1154
rect 6072 -1188 6106 -1154
rect 6140 -1188 6174 -1154
rect 6208 -1188 6242 -1154
rect 6276 -1188 6310 -1154
rect 6344 -1188 6378 -1154
rect 6412 -1188 6446 -1154
rect 6480 -1188 6514 -1154
rect 6548 -1188 6582 -1154
rect 6616 -1188 6650 -1154
rect 6684 -1188 6718 -1154
rect 6752 -1188 6786 -1154
rect 6820 -1188 6854 -1154
rect 6888 -1188 6922 -1154
rect 6956 -1188 6990 -1154
rect 7024 -1188 7058 -1154
rect 7092 -1188 7126 -1154
rect 7160 -1188 7194 -1154
rect 7228 -1188 7262 -1154
rect 7296 -1188 7330 -1154
rect 7364 -1188 7398 -1154
rect 7432 -1188 7466 -1154
rect 7500 -1188 7534 -1154
rect 7568 -1188 7602 -1154
rect 7636 -1188 7670 -1154
rect 7704 -1188 7738 -1154
rect 7772 -1188 7806 -1154
rect 7840 -1188 7874 -1154
rect 7908 -1188 7976 -1154
rect 5617 -1222 5651 -1188
rect 5617 -1290 5651 -1256
rect 7942 -1262 7976 -1188
rect 5617 -1358 5651 -1324
rect 5617 -1426 5651 -1392
rect 5617 -1494 5651 -1460
rect 5617 -1562 5651 -1528
rect 5617 -1724 5651 -1596
rect 5617 -1792 5651 -1758
rect 5617 -1860 5651 -1826
rect 7942 -1330 7976 -1296
rect 7942 -1398 7976 -1364
rect 7942 -1466 7976 -1432
rect 7942 -1534 7976 -1500
rect 7942 -1602 7976 -1568
rect 7942 -1670 7976 -1636
rect 7942 -1738 7976 -1704
rect 7942 -1806 7976 -1772
rect 7942 -1874 7976 -1840
rect 5617 -1928 5651 -1894
rect 5617 -2010 5651 -1962
rect 7942 -1942 7976 -1908
rect 7942 -2010 7976 -1976
rect 5617 -2044 5685 -2010
rect 5719 -2044 5753 -2010
rect 5787 -2044 5821 -2010
rect 5855 -2044 5889 -2010
rect 5923 -2044 5957 -2010
rect 5991 -2044 6025 -2010
rect 6059 -2044 6093 -2010
rect 6127 -2044 6161 -2010
rect 6195 -2044 6229 -2010
rect 6263 -2044 6297 -2010
rect 6331 -2044 6365 -2010
rect 6399 -2044 6433 -2010
rect 6467 -2044 6501 -2010
rect 6535 -2044 6569 -2010
rect 6603 -2044 6637 -2010
rect 6671 -2044 6705 -2010
rect 6739 -2044 6773 -2010
rect 6807 -2044 6841 -2010
rect 6875 -2044 6909 -2010
rect 6943 -2044 6977 -2010
rect 7011 -2044 7045 -2010
rect 7079 -2044 7113 -2010
rect 7147 -2044 7181 -2010
rect 7215 -2044 7249 -2010
rect 7283 -2044 7317 -2010
rect 7351 -2044 7385 -2010
rect 7419 -2044 7453 -2010
rect 7487 -2044 7521 -2010
rect 7555 -2044 7589 -2010
rect 7623 -2044 7657 -2010
rect 7691 -2044 7725 -2010
rect 7759 -2044 7793 -2010
rect 7827 -2044 7861 -2010
rect 7895 -2044 7976 -2010
<< mvpsubdiffcont >>
rect 458 1317 492 1351
rect 526 1317 560 1351
rect 594 1317 628 1351
rect 662 1317 696 1351
rect 730 1317 764 1351
rect 798 1317 832 1351
rect 866 1317 900 1351
rect 934 1317 968 1351
rect 1002 1317 1036 1351
rect 1131 1317 1165 1351
rect 1199 1317 1233 1351
rect 1267 1317 1301 1351
rect 1335 1317 1369 1351
rect 1403 1317 1437 1351
rect 1471 1317 1505 1351
rect 1539 1317 1573 1351
rect 1607 1317 1641 1351
rect 360 1252 394 1286
rect 360 1184 394 1218
rect 360 1116 394 1150
rect 360 1048 394 1082
rect 360 980 394 1014
rect 360 912 394 946
rect 360 844 394 878
rect 360 776 394 810
rect 360 708 394 742
rect 360 640 394 674
rect 360 572 394 606
rect 1672 1206 1706 1240
rect 1672 1138 1706 1172
rect 1672 1070 1706 1104
rect 1672 1002 1706 1036
rect 1672 934 1706 968
rect 1672 866 1706 900
rect 1672 798 1706 832
rect 1672 730 1706 764
rect 1672 662 1706 696
rect 1672 594 1706 628
rect 360 504 394 538
rect 1672 526 1706 560
rect 360 436 394 470
rect 1672 458 1706 492
rect 1672 390 1706 424
rect 425 325 459 359
rect 493 325 527 359
rect 561 325 595 359
rect 629 325 663 359
rect 697 325 731 359
rect 765 325 799 359
rect 833 325 867 359
rect 901 325 935 359
rect 969 325 1003 359
rect 1037 325 1071 359
rect 1105 325 1139 359
rect 1173 325 1207 359
rect 1241 325 1275 359
rect 1309 325 1343 359
rect 1377 325 1411 359
rect 1445 325 1479 359
rect 1513 325 1547 359
rect 1581 325 1615 359
rect 2287 1343 2321 1377
rect 2355 1343 2389 1377
rect 2423 1343 2457 1377
rect 2491 1343 2525 1377
rect 2559 1343 2593 1377
rect 2627 1343 2661 1377
rect 2695 1343 2729 1377
rect 2763 1343 2797 1377
rect 2831 1343 2865 1377
rect 2899 1343 2933 1377
rect 2967 1343 3001 1377
rect 3035 1343 3069 1377
rect 3103 1343 3137 1377
rect 3171 1343 3205 1377
rect 3239 1343 3273 1377
rect 3307 1343 3341 1377
rect 3375 1343 3409 1377
rect 3443 1343 3477 1377
rect 3511 1343 3545 1377
rect 3579 1343 3613 1377
rect 3647 1343 3681 1377
rect 3715 1343 3749 1377
rect 3783 1343 3817 1377
rect 3851 1343 3885 1377
rect 3919 1343 3953 1377
rect 3987 1343 4021 1377
rect 4055 1343 4089 1377
rect 4123 1343 4157 1377
rect 4191 1343 4225 1377
rect 4259 1343 4293 1377
rect 4327 1343 4361 1377
rect 4395 1343 4429 1377
rect 4558 1343 4592 1377
rect 4626 1343 4660 1377
rect 4694 1343 4728 1377
rect 4762 1343 4796 1377
rect 4830 1343 4864 1377
rect 4898 1343 4932 1377
rect 4966 1343 5000 1377
rect 5034 1343 5068 1377
rect 5102 1343 5136 1377
rect 5170 1343 5204 1377
rect 5238 1343 5272 1377
rect 5306 1343 5340 1377
rect 5374 1343 5408 1377
rect 5442 1343 5476 1377
rect 5510 1343 5544 1377
rect 5578 1343 5612 1377
rect 5646 1343 5680 1377
rect 5714 1343 5748 1377
rect 5782 1343 5816 1377
rect 5850 1343 5884 1377
rect 5918 1343 5952 1377
rect 5986 1343 6020 1377
rect 6054 1343 6088 1377
rect 6122 1343 6156 1377
rect 6190 1343 6224 1377
rect 6258 1343 6292 1377
rect 6326 1343 6360 1377
rect 6394 1343 6428 1377
rect 6462 1343 6496 1377
rect 6530 1343 6564 1377
rect 6598 1343 6632 1377
rect 2195 1278 2229 1312
rect 6663 1274 6697 1308
rect 2195 1210 2229 1244
rect 2195 1142 2229 1176
rect 2195 1074 2229 1108
rect 2195 1006 2229 1040
rect 2195 938 2229 972
rect 2195 870 2229 904
rect 2195 802 2229 836
rect 2195 734 2229 768
rect 2195 666 2229 700
rect 2195 598 2229 632
rect 2195 530 2229 564
rect 2195 462 2229 496
rect 6663 1206 6697 1240
rect 6663 1138 6697 1172
rect 6663 1070 6697 1104
rect 6663 1002 6697 1036
rect 6663 934 6697 968
rect 6663 866 6697 900
rect 6663 798 6697 832
rect 6663 730 6697 764
rect 6663 662 6697 696
rect 6663 594 6697 628
rect 6663 526 6697 560
rect 6663 458 6697 492
rect 2195 394 2229 428
rect 6663 390 6697 424
rect 2260 325 2294 359
rect 2328 325 2362 359
rect 2396 325 2430 359
rect 2464 325 2498 359
rect 2532 325 2566 359
rect 2600 325 2634 359
rect 2668 325 2702 359
rect 2736 325 2770 359
rect 2804 325 2838 359
rect 2872 325 2906 359
rect 2940 325 2974 359
rect 3008 325 3042 359
rect 3076 325 3110 359
rect 3144 325 3178 359
rect 3212 325 3246 359
rect 3280 325 3314 359
rect 3348 325 3382 359
rect 3416 325 3450 359
rect 3484 325 3518 359
rect 3552 325 3586 359
rect 3620 325 3654 359
rect 3688 325 3722 359
rect 3756 325 3790 359
rect 3824 325 3858 359
rect 3892 325 3926 359
rect 3960 325 3994 359
rect 4028 325 4062 359
rect 4096 325 4130 359
rect 4164 325 4198 359
rect 4232 325 4266 359
rect 4300 325 4334 359
rect 4368 325 4402 359
rect 4436 325 4470 359
rect 4504 325 4538 359
rect 4572 325 4606 359
rect 4640 325 4674 359
rect 4708 325 4742 359
rect 4776 325 4810 359
rect 4844 325 4878 359
rect 4912 325 4946 359
rect 4980 325 5014 359
rect 5048 325 5082 359
rect 5116 325 5150 359
rect 5184 325 5218 359
rect 5252 325 5286 359
rect 5320 325 5354 359
rect 5388 325 5422 359
rect 5456 325 5490 359
rect 5524 325 5558 359
rect 5592 325 5626 359
rect 5660 325 5694 359
rect 5728 325 5762 359
rect 5796 325 5830 359
rect 5864 325 5898 359
rect 5932 325 5966 359
rect 6000 325 6034 359
rect 6068 325 6102 359
rect 6136 325 6170 359
rect 6204 325 6238 359
rect 6272 325 6306 359
rect 6340 325 6374 359
rect 6408 325 6442 359
rect 6476 325 6510 359
rect 6544 325 6578 359
rect 7264 1343 7298 1377
rect 7332 1343 7366 1377
rect 7400 1343 7434 1377
rect 7468 1343 7502 1377
rect 7536 1343 7570 1377
rect 7604 1343 7638 1377
rect 7672 1343 7706 1377
rect 7740 1343 7774 1377
rect 7808 1343 7842 1377
rect 7876 1343 7910 1377
rect 7944 1343 7978 1377
rect 8012 1343 8046 1377
rect 8080 1343 8114 1377
rect 8148 1343 8182 1377
rect 8216 1343 8250 1377
rect 8284 1343 8318 1377
rect 8352 1343 8386 1377
rect 8420 1343 8454 1377
rect 8488 1343 8522 1377
rect 8556 1343 8590 1377
rect 8624 1343 8658 1377
rect 8692 1343 8726 1377
rect 8760 1343 8794 1377
rect 8828 1343 8862 1377
rect 8896 1343 8930 1377
rect 8964 1343 8998 1377
rect 9032 1343 9066 1377
rect 9100 1343 9134 1377
rect 9168 1343 9202 1377
rect 9236 1343 9270 1377
rect 9304 1343 9338 1377
rect 9372 1343 9406 1377
rect 9500 1343 9534 1377
rect 9568 1343 9602 1377
rect 9636 1343 9670 1377
rect 9704 1343 9738 1377
rect 9772 1343 9806 1377
rect 9840 1343 9874 1377
rect 9908 1343 9942 1377
rect 9976 1343 10010 1377
rect 10044 1343 10078 1377
rect 10112 1343 10146 1377
rect 10180 1343 10214 1377
rect 10248 1343 10282 1377
rect 10316 1343 10350 1377
rect 10384 1343 10418 1377
rect 10452 1343 10486 1377
rect 10520 1343 10554 1377
rect 10588 1343 10622 1377
rect 10656 1343 10690 1377
rect 10724 1343 10758 1377
rect 10792 1343 10826 1377
rect 10860 1343 10894 1377
rect 10928 1343 10962 1377
rect 10996 1343 11030 1377
rect 11064 1343 11098 1377
rect 11132 1343 11166 1377
rect 11200 1343 11234 1377
rect 11268 1343 11302 1377
rect 11336 1343 11370 1377
rect 11404 1343 11438 1377
rect 11472 1343 11506 1377
rect 11540 1343 11574 1377
rect 11608 1343 11642 1377
rect 7199 1274 7233 1308
rect 11681 1278 11715 1312
rect 7199 1206 7233 1240
rect 7199 1138 7233 1172
rect 7199 1070 7233 1104
rect 7199 1002 7233 1036
rect 7199 934 7233 968
rect 7199 866 7233 900
rect 7199 798 7233 832
rect 7199 730 7233 764
rect 7199 662 7233 696
rect 7199 594 7233 628
rect 7199 526 7233 560
rect 7199 458 7233 492
rect 11681 1210 11715 1244
rect 11681 1142 11715 1176
rect 11681 1074 11715 1108
rect 11681 1006 11715 1040
rect 11681 938 11715 972
rect 11681 870 11715 904
rect 11681 802 11715 836
rect 11681 734 11715 768
rect 11681 666 11715 700
rect 11681 598 11715 632
rect 11681 530 11715 564
rect 11681 462 11715 496
rect 7199 390 7233 424
rect 11681 394 11715 428
rect 7264 325 7298 359
rect 7332 325 7366 359
rect 7400 325 7434 359
rect 7468 325 7502 359
rect 7536 325 7570 359
rect 7604 325 7638 359
rect 7672 325 7706 359
rect 7740 325 7774 359
rect 7808 325 7842 359
rect 7876 325 7910 359
rect 7944 325 7978 359
rect 8012 325 8046 359
rect 8080 325 8114 359
rect 8148 325 8182 359
rect 8216 325 8250 359
rect 8284 325 8318 359
rect 8352 325 8386 359
rect 8420 325 8454 359
rect 8488 325 8522 359
rect 8556 325 8590 359
rect 8624 325 8658 359
rect 8692 325 8726 359
rect 8760 325 8794 359
rect 8828 325 8862 359
rect 8896 325 8930 359
rect 8964 325 8998 359
rect 9032 325 9066 359
rect 9100 325 9134 359
rect 9168 325 9202 359
rect 9236 325 9270 359
rect 9304 325 9338 359
rect 9372 325 9406 359
rect 9440 325 9474 359
rect 9508 325 9542 359
rect 9576 325 9610 359
rect 9644 325 9678 359
rect 9712 325 9746 359
rect 9780 325 9814 359
rect 9848 325 9882 359
rect 9916 325 9950 359
rect 9984 325 10018 359
rect 10052 325 10086 359
rect 10120 325 10154 359
rect 10188 325 10222 359
rect 10256 325 10290 359
rect 10324 325 10358 359
rect 10392 325 10426 359
rect 10460 325 10494 359
rect 10528 325 10562 359
rect 10596 325 10630 359
rect 10664 325 10698 359
rect 10732 325 10766 359
rect 10800 325 10834 359
rect 10868 325 10902 359
rect 10936 325 10970 359
rect 11004 325 11038 359
rect 11072 325 11106 359
rect 11140 325 11174 359
rect 11208 325 11242 359
rect 11276 325 11310 359
rect 11344 325 11378 359
rect 11412 325 11446 359
rect 11480 325 11514 359
rect 11548 325 11582 359
rect 11616 325 11650 359
<< mvnsubdiffcont >>
rect 63 135 165 1461
rect 138 67 172 101
rect 206 67 1872 169
rect 1906 135 2008 1461
rect 6884 260 6986 1450
rect 2035 67 2069 101
rect 2103 67 4653 169
rect 7020 135 7054 169
rect 7089 135 7123 169
rect 7158 135 7192 169
rect 7227 135 7261 169
rect 7296 135 7330 169
rect 7365 135 7399 169
rect 7434 135 7468 169
rect 7503 135 7537 169
rect 7572 135 7606 169
rect 7641 135 7675 169
rect 7710 135 7744 169
rect 7779 135 7813 169
rect 7848 135 7882 169
rect 7917 135 7951 169
rect 7986 135 8020 169
rect 8055 135 8089 169
rect 8124 135 8158 169
rect 8193 135 8227 169
rect 8262 135 8296 169
rect 8331 135 8365 169
rect 8400 135 8434 169
rect 8469 135 8503 169
rect 8538 135 8572 169
rect 8607 135 8641 169
rect 8676 135 8710 169
rect 8745 135 8779 169
rect 8814 135 8848 169
rect 8883 135 8917 169
rect 7020 67 7054 101
rect 7089 67 7123 101
rect 7158 67 7192 101
rect 7227 67 7261 101
rect 7296 67 7330 101
rect 7365 67 7399 101
rect 7434 67 7468 101
rect 7503 67 7537 101
rect 7572 67 7606 101
rect 7641 67 7675 101
rect 7710 67 7744 101
rect 7779 67 7813 101
rect 7848 67 7882 101
rect 7917 67 7951 101
rect 7986 67 8020 101
rect 8055 67 8089 101
rect 8124 67 8158 101
rect 8193 67 8227 101
rect 8262 67 8296 101
rect 8331 67 8365 101
rect 8400 67 8434 101
rect 8469 67 8503 101
rect 8538 67 8572 101
rect 8607 67 8641 101
rect 8676 67 8710 101
rect 8745 67 8779 101
rect 8814 67 8848 101
rect 8883 67 8917 101
rect 8952 67 11842 169
rect 5698 -1188 5732 -1154
rect 5766 -1188 5800 -1154
rect 5834 -1188 5868 -1154
rect 5902 -1188 5936 -1154
rect 5970 -1188 6004 -1154
rect 6038 -1188 6072 -1154
rect 6106 -1188 6140 -1154
rect 6174 -1188 6208 -1154
rect 6242 -1188 6276 -1154
rect 6310 -1188 6344 -1154
rect 6378 -1188 6412 -1154
rect 6446 -1188 6480 -1154
rect 6514 -1188 6548 -1154
rect 6582 -1188 6616 -1154
rect 6650 -1188 6684 -1154
rect 6718 -1188 6752 -1154
rect 6786 -1188 6820 -1154
rect 6854 -1188 6888 -1154
rect 6922 -1188 6956 -1154
rect 6990 -1188 7024 -1154
rect 7058 -1188 7092 -1154
rect 7126 -1188 7160 -1154
rect 7194 -1188 7228 -1154
rect 7262 -1188 7296 -1154
rect 7330 -1188 7364 -1154
rect 7398 -1188 7432 -1154
rect 7466 -1188 7500 -1154
rect 7534 -1188 7568 -1154
rect 7602 -1188 7636 -1154
rect 7670 -1188 7704 -1154
rect 7738 -1188 7772 -1154
rect 7806 -1188 7840 -1154
rect 7874 -1188 7908 -1154
rect 5617 -1256 5651 -1222
rect 5617 -1324 5651 -1290
rect 7942 -1296 7976 -1262
rect 5617 -1392 5651 -1358
rect 5617 -1460 5651 -1426
rect 5617 -1528 5651 -1494
rect 5617 -1596 5651 -1562
rect 5617 -1758 5651 -1724
rect 5617 -1826 5651 -1792
rect 5617 -1894 5651 -1860
rect 7942 -1364 7976 -1330
rect 7942 -1432 7976 -1398
rect 7942 -1500 7976 -1466
rect 7942 -1568 7976 -1534
rect 7942 -1636 7976 -1602
rect 7942 -1704 7976 -1670
rect 7942 -1772 7976 -1738
rect 7942 -1840 7976 -1806
rect 5617 -1962 5651 -1928
rect 7942 -1908 7976 -1874
rect 7942 -1976 7976 -1942
rect 5685 -2044 5719 -2010
rect 5753 -2044 5787 -2010
rect 5821 -2044 5855 -2010
rect 5889 -2044 5923 -2010
rect 5957 -2044 5991 -2010
rect 6025 -2044 6059 -2010
rect 6093 -2044 6127 -2010
rect 6161 -2044 6195 -2010
rect 6229 -2044 6263 -2010
rect 6297 -2044 6331 -2010
rect 6365 -2044 6399 -2010
rect 6433 -2044 6467 -2010
rect 6501 -2044 6535 -2010
rect 6569 -2044 6603 -2010
rect 6637 -2044 6671 -2010
rect 6705 -2044 6739 -2010
rect 6773 -2044 6807 -2010
rect 6841 -2044 6875 -2010
rect 6909 -2044 6943 -2010
rect 6977 -2044 7011 -2010
rect 7045 -2044 7079 -2010
rect 7113 -2044 7147 -2010
rect 7181 -2044 7215 -2010
rect 7249 -2044 7283 -2010
rect 7317 -2044 7351 -2010
rect 7385 -2044 7419 -2010
rect 7453 -2044 7487 -2010
rect 7521 -2044 7555 -2010
rect 7589 -2044 7623 -2010
rect 7657 -2044 7691 -2010
rect 7725 -2044 7759 -2010
rect 7793 -2044 7827 -2010
rect 7861 -2044 7895 -2010
<< poly >>
rect -506 686 -106 688
rect 460 1230 526 1246
rect 460 1196 476 1230
rect 510 1196 526 1230
rect 460 1187 526 1196
rect 460 1160 558 1187
rect 460 1126 476 1160
rect 510 1126 558 1160
rect 460 1090 558 1126
rect 460 1056 476 1090
rect 510 1087 558 1090
rect 1558 1087 1590 1187
rect 510 1056 526 1087
rect 460 1031 526 1056
rect 460 1020 558 1031
rect 460 986 476 1020
rect 510 986 558 1020
rect 460 950 558 986
rect 460 916 476 950
rect 510 931 558 950
rect 1558 931 1590 1031
rect 510 916 526 931
rect 460 880 526 916
rect 460 846 476 880
rect 510 846 526 880
rect 460 810 526 846
rect 460 776 476 810
rect 510 776 526 810
rect 460 745 526 776
rect 460 740 558 745
rect 460 706 476 740
rect 510 706 558 740
rect 460 669 558 706
rect 460 635 476 669
rect 510 645 558 669
rect 1558 645 1590 745
rect 510 635 526 645
rect 460 598 526 635
rect 460 564 476 598
rect 510 589 526 598
rect 510 564 558 589
rect 460 548 558 564
rect 526 489 558 548
rect 1558 489 1590 589
rect 2295 1197 2393 1213
rect 2295 1163 2311 1197
rect 2345 1163 2393 1197
rect 2295 1123 2393 1163
rect 2295 1089 2311 1123
rect 2345 1113 2393 1123
rect 4393 1113 4425 1213
rect 4467 1113 4499 1213
rect 6499 1197 6597 1213
rect 6499 1163 6547 1197
rect 6581 1163 6597 1197
rect 6499 1123 6597 1163
rect 6499 1113 6547 1123
rect 2345 1089 2361 1113
rect 2295 1057 2361 1089
rect 6531 1089 6547 1113
rect 6581 1089 6597 1123
rect 6531 1057 6597 1089
rect 2295 1049 2393 1057
rect 2295 1015 2311 1049
rect 2345 1015 2393 1049
rect 2295 974 2393 1015
rect 2295 940 2311 974
rect 2345 957 2393 974
rect 4393 957 4425 1057
rect 4467 957 4499 1057
rect 6499 1049 6597 1057
rect 6499 1015 6547 1049
rect 6581 1015 6597 1049
rect 6499 974 6597 1015
rect 6499 957 6547 974
rect 2345 940 2361 957
rect 2295 901 2361 940
rect 6531 940 6547 957
rect 6581 940 6597 974
rect 6531 901 6597 940
rect 2295 899 2393 901
rect 2295 865 2311 899
rect 2345 865 2393 899
rect 2295 824 2393 865
rect 2295 790 2311 824
rect 2345 801 2393 824
rect 4393 801 4425 901
rect 4467 801 4499 901
rect 6499 899 6597 901
rect 6499 865 6547 899
rect 6581 865 6597 899
rect 6499 824 6597 865
rect 6499 801 6547 824
rect 2345 790 2361 801
rect 2295 749 2361 790
rect 2295 715 2311 749
rect 2345 745 2361 749
rect 6531 790 6547 801
rect 6581 790 6597 824
rect 6531 749 6597 790
rect 6531 745 6547 749
rect 2345 715 2393 745
rect 2295 674 2393 715
rect 2295 640 2311 674
rect 2345 645 2393 674
rect 4393 645 4425 745
rect 4467 645 4499 745
rect 6499 715 6547 745
rect 6581 715 6597 749
rect 6499 674 6597 715
rect 6499 645 6547 674
rect 2345 640 2361 645
rect 2295 599 2361 640
rect 2295 565 2311 599
rect 2345 589 2361 599
rect 6531 640 6547 645
rect 6581 640 6597 674
rect 6531 599 6597 640
rect 6531 589 6547 599
rect 2345 565 2393 589
rect 2295 549 2393 565
rect 2361 489 2393 549
rect 4393 489 4425 589
rect 4467 489 4499 589
rect 6499 565 6547 589
rect 6581 565 6597 599
rect 6499 549 6597 565
rect 6499 489 6531 549
rect 7314 1197 7412 1213
rect 7314 1163 7330 1197
rect 7364 1163 7412 1197
rect 7314 1123 7412 1163
rect 7314 1089 7330 1123
rect 7364 1113 7412 1123
rect 9412 1113 9444 1213
rect 9486 1113 9518 1213
rect 11518 1197 11615 1213
rect 11518 1163 11565 1197
rect 11599 1163 11615 1197
rect 11518 1123 11615 1163
rect 11518 1113 11565 1123
rect 7364 1089 7380 1113
rect 7314 1057 7380 1089
rect 11549 1089 11565 1113
rect 11599 1089 11615 1123
rect 11549 1057 11615 1089
rect 7314 1050 7412 1057
rect 7314 1016 7330 1050
rect 7364 1016 7412 1050
rect 7314 977 7412 1016
rect 7314 943 7330 977
rect 7364 957 7412 977
rect 9412 957 9444 1057
rect 9486 957 9518 1057
rect 11518 1050 11615 1057
rect 11518 1016 11565 1050
rect 11599 1016 11615 1050
rect 11518 977 11615 1016
rect 11518 957 11565 977
rect 7364 943 7380 957
rect 7314 904 7380 943
rect 7314 870 7330 904
rect 7364 901 7380 904
rect 11549 943 11565 957
rect 11599 943 11615 977
rect 11549 904 11615 943
rect 11549 901 11565 904
rect 7364 870 7412 901
rect 7314 831 7412 870
rect 7314 797 7330 831
rect 7364 801 7412 831
rect 9412 801 9444 901
rect 9486 801 9518 901
rect 11518 870 11565 901
rect 11599 870 11615 904
rect 11518 831 11615 870
rect 11518 801 11565 831
rect 7364 797 7380 801
rect 7314 758 7380 797
rect 7314 724 7330 758
rect 7364 745 7380 758
rect 11549 797 11565 801
rect 11599 797 11615 831
rect 11549 758 11615 797
rect 11549 745 11565 758
rect 7364 724 7412 745
rect 7314 685 7412 724
rect 7314 651 7330 685
rect 7364 651 7412 685
rect 7314 645 7412 651
rect 9412 645 9444 745
rect 9486 645 9518 745
rect 11518 724 11565 745
rect 11599 724 11615 758
rect 11518 685 11615 724
rect 11518 651 11565 685
rect 11599 651 11615 685
rect 11518 645 11615 651
rect 7314 612 7380 645
rect 7314 578 7330 612
rect 7364 589 7380 612
rect 11549 612 11615 645
rect 11549 589 11565 612
rect 7364 578 7412 589
rect 7314 539 7412 578
rect 7314 505 7330 539
rect 7364 505 7412 539
rect 7314 489 7412 505
rect 9412 489 9444 589
rect 9486 489 9518 589
rect 11518 578 11565 589
rect 11599 578 11615 612
rect 11518 539 11615 578
rect 11518 505 11565 539
rect 11599 505 11615 539
rect 11518 489 11615 505
rect 5718 -1331 5816 -1315
rect 5718 -1365 5734 -1331
rect 5768 -1365 5816 -1331
rect 5718 -1402 5816 -1365
rect 5718 -1436 5734 -1402
rect 5768 -1415 5816 -1402
rect 7816 -1415 7848 -1315
rect 5768 -1436 5784 -1415
rect 5718 -1471 5784 -1436
rect 5718 -1473 5816 -1471
rect 5718 -1507 5734 -1473
rect 5768 -1507 5816 -1473
rect 5718 -1545 5816 -1507
rect 5718 -1579 5734 -1545
rect 5768 -1571 5816 -1545
rect 7816 -1571 7848 -1471
rect 5768 -1579 5784 -1571
rect 5718 -1617 5784 -1579
rect 5718 -1651 5734 -1617
rect 5768 -1627 5784 -1617
rect 5768 -1651 5816 -1627
rect 5718 -1689 5816 -1651
rect 5718 -1723 5734 -1689
rect 5768 -1723 5816 -1689
rect 5718 -1727 5816 -1723
rect 7816 -1727 7848 -1627
rect 5718 -1761 5784 -1727
rect 5718 -1795 5734 -1761
rect 5768 -1783 5784 -1761
rect 5768 -1795 5816 -1783
rect 5718 -1833 5816 -1795
rect 5718 -1867 5734 -1833
rect 5768 -1867 5816 -1833
rect 5718 -1883 5816 -1867
rect 7816 -1883 7848 -1783
<< polycont >>
rect 476 1196 510 1230
rect 476 1126 510 1160
rect 476 1056 510 1090
rect 476 986 510 1020
rect 476 916 510 950
rect 476 846 510 880
rect 476 776 510 810
rect 476 706 510 740
rect 476 635 510 669
rect 476 564 510 598
rect 2311 1163 2345 1197
rect 2311 1089 2345 1123
rect 6547 1163 6581 1197
rect 6547 1089 6581 1123
rect 2311 1015 2345 1049
rect 2311 940 2345 974
rect 6547 1015 6581 1049
rect 6547 940 6581 974
rect 2311 865 2345 899
rect 2311 790 2345 824
rect 6547 865 6581 899
rect 2311 715 2345 749
rect 6547 790 6581 824
rect 2311 640 2345 674
rect 6547 715 6581 749
rect 2311 565 2345 599
rect 6547 640 6581 674
rect 6547 565 6581 599
rect 7330 1163 7364 1197
rect 7330 1089 7364 1123
rect 11565 1163 11599 1197
rect 11565 1089 11599 1123
rect 7330 1016 7364 1050
rect 7330 943 7364 977
rect 11565 1016 11599 1050
rect 7330 870 7364 904
rect 11565 943 11599 977
rect 7330 797 7364 831
rect 11565 870 11599 904
rect 7330 724 7364 758
rect 11565 797 11599 831
rect 7330 651 7364 685
rect 11565 724 11599 758
rect 11565 651 11599 685
rect 7330 578 7364 612
rect 7330 505 7364 539
rect 11565 578 11599 612
rect 11565 505 11599 539
rect 5734 -1365 5768 -1331
rect 5734 -1436 5768 -1402
rect 5734 -1507 5768 -1473
rect 5734 -1579 5768 -1545
rect 5734 -1651 5768 -1617
rect 5734 -1723 5768 -1689
rect 5734 -1795 5768 -1761
rect 5734 -1867 5768 -1833
<< locali >>
rect 63 1534 6986 1636
rect -462 1460 -409 1494
rect -375 1460 -322 1494
rect -288 1460 -236 1494
rect -202 1460 -150 1494
rect -496 1384 -116 1460
rect 63 1461 165 1534
rect 1906 1466 2008 1534
rect -462 1350 -409 1384
rect -375 1350 -322 1384
rect -288 1350 -236 1384
rect -202 1350 -150 1384
rect 55 1408 63 1446
rect 1898 1461 2016 1466
rect 165 1408 173 1446
rect 1898 1434 1906 1461
rect 2008 1434 2016 1461
rect 55 1374 61 1408
rect 167 1374 173 1408
rect 55 1335 63 1374
rect 165 1335 173 1374
rect 55 1301 61 1335
rect 167 1301 173 1335
rect 55 1262 63 1301
rect 165 1262 173 1301
rect 55 1228 61 1262
rect 167 1228 173 1262
rect 55 1189 63 1228
rect 165 1189 173 1228
rect 55 1155 61 1189
rect 167 1155 173 1189
rect 55 1116 63 1155
rect 165 1116 173 1155
rect 55 1082 61 1116
rect 167 1082 173 1116
rect 55 1043 63 1082
rect 165 1043 173 1082
rect 55 1009 61 1043
rect 167 1009 173 1043
rect 55 970 63 1009
rect 165 970 173 1009
rect 55 936 61 970
rect 167 936 173 970
rect 55 897 63 936
rect 165 897 173 936
rect 55 863 61 897
rect 167 863 173 897
rect 55 824 63 863
rect 165 824 173 863
rect 55 790 61 824
rect 167 790 173 824
rect -463 726 -410 760
rect -376 726 -323 760
rect -289 726 -236 760
rect -202 726 -150 760
rect -497 682 -116 726
rect -463 648 -410 682
rect -376 648 -323 682
rect -289 648 -236 682
rect -202 648 -150 682
rect -497 604 -116 648
rect -463 570 -410 604
rect -376 570 -323 604
rect -289 570 -236 604
rect -202 570 -150 604
rect 55 751 63 790
rect 165 751 173 790
rect 55 717 61 751
rect 167 717 173 751
rect 55 678 63 717
rect 165 678 173 717
rect 55 644 61 678
rect 167 644 173 678
rect 55 605 63 644
rect 165 605 173 644
rect 55 571 61 605
rect 167 571 173 605
rect 55 532 63 571
rect 165 532 173 571
rect 55 498 61 532
rect 167 498 173 532
rect 55 459 63 498
rect 165 459 173 498
rect 55 137 61 459
rect 167 177 173 459
rect 318 1426 1748 1432
rect 318 1392 402 1426
rect 436 1392 480 1426
rect 514 1392 558 1426
rect 592 1392 636 1426
rect 670 1392 714 1426
rect 748 1392 792 1426
rect 826 1392 870 1426
rect 904 1392 949 1426
rect 983 1392 1059 1426
rect 318 1354 1059 1392
rect 318 1320 324 1354
rect 358 1320 396 1354
rect 430 1351 480 1354
rect 514 1351 558 1354
rect 592 1351 636 1354
rect 670 1351 714 1354
rect 748 1351 792 1354
rect 826 1351 870 1354
rect 904 1351 949 1354
rect 983 1351 1059 1354
rect 1597 1392 1636 1426
rect 1670 1392 1748 1426
rect 1597 1354 1748 1392
rect 1597 1351 1636 1354
rect 430 1320 458 1351
rect 514 1320 526 1351
rect 592 1320 594 1351
rect 318 1317 458 1320
rect 492 1317 526 1320
rect 560 1317 594 1320
rect 628 1320 636 1351
rect 696 1320 714 1351
rect 764 1320 792 1351
rect 628 1317 662 1320
rect 696 1317 730 1320
rect 764 1317 798 1320
rect 832 1317 866 1351
rect 904 1320 934 1351
rect 983 1320 1002 1351
rect 900 1317 934 1320
rect 968 1317 1002 1320
rect 1036 1320 1059 1351
rect 1597 1320 1607 1351
rect 1670 1350 1748 1354
rect 1670 1320 1708 1350
rect 1036 1317 1131 1320
rect 1165 1317 1199 1320
rect 1233 1317 1267 1320
rect 1301 1317 1335 1320
rect 1369 1317 1403 1320
rect 1437 1317 1471 1320
rect 1505 1317 1539 1320
rect 1573 1317 1607 1320
rect 1641 1317 1708 1320
rect 318 1316 1708 1317
rect 1742 1316 1748 1350
rect 318 1314 1748 1316
rect 318 1286 436 1314
rect 318 1277 360 1286
rect 318 1243 324 1277
rect 358 1252 360 1277
rect 394 1277 436 1286
rect 394 1252 396 1277
rect 358 1243 396 1252
rect 430 1243 436 1277
rect 1630 1274 1748 1314
rect 318 1218 436 1243
rect 318 1200 360 1218
rect 318 1166 324 1200
rect 358 1184 360 1200
rect 394 1200 436 1218
rect 394 1184 396 1200
rect 358 1166 396 1184
rect 430 1166 436 1200
rect 318 1150 436 1166
rect 318 1123 360 1150
rect 318 1089 324 1123
rect 358 1116 360 1123
rect 394 1123 436 1150
rect 394 1116 396 1123
rect 358 1089 396 1116
rect 430 1089 436 1123
rect 318 1082 436 1089
rect 318 1048 360 1082
rect 394 1048 436 1082
rect 318 1046 436 1048
rect 318 1012 324 1046
rect 358 1014 396 1046
rect 358 1012 360 1014
rect 318 980 360 1012
rect 394 1012 396 1014
rect 430 1012 436 1046
rect 394 980 436 1012
rect 318 969 436 980
rect 318 935 324 969
rect 358 946 396 969
rect 358 935 360 946
rect 318 912 360 935
rect 394 935 396 946
rect 430 935 436 969
rect 394 912 436 935
rect 318 892 436 912
rect 318 858 324 892
rect 358 878 396 892
rect 358 858 360 878
rect 318 844 360 858
rect 394 858 396 878
rect 430 858 436 892
rect 394 844 436 858
rect 318 816 436 844
rect 318 782 324 816
rect 358 810 396 816
rect 358 782 360 810
rect 318 776 360 782
rect 394 782 396 810
rect 430 782 436 816
rect 394 776 436 782
rect 318 742 436 776
rect 318 740 360 742
rect 318 706 324 740
rect 358 708 360 740
rect 394 740 436 742
rect 394 708 396 740
rect 358 706 396 708
rect 430 706 436 740
rect 318 674 436 706
rect 318 664 360 674
rect 318 630 324 664
rect 358 640 360 664
rect 394 664 436 674
rect 394 640 396 664
rect 358 630 396 640
rect 430 630 436 664
rect 318 606 436 630
rect 318 588 360 606
rect 318 554 324 588
rect 358 572 360 588
rect 394 588 436 606
rect 394 572 396 588
rect 358 554 396 572
rect 430 554 436 588
rect 318 538 436 554
rect 318 512 360 538
rect 318 478 324 512
rect 358 504 360 512
rect 394 512 436 538
rect 394 504 396 512
rect 358 478 396 504
rect 430 478 436 512
rect 476 1230 510 1246
rect 1630 1240 1636 1274
rect 1670 1240 1708 1274
rect 1742 1240 1748 1274
rect 600 1232 641 1235
rect 675 1232 716 1235
rect 750 1232 791 1235
rect 825 1232 866 1235
rect 900 1232 940 1235
rect 974 1232 1014 1235
rect 1048 1232 1088 1235
rect 1122 1232 1162 1235
rect 1196 1232 1236 1235
rect 1270 1232 1310 1235
rect 1344 1232 1384 1235
rect 1418 1232 1458 1235
rect 554 1201 566 1232
rect 554 1198 570 1201
rect 604 1198 638 1232
rect 675 1201 706 1232
rect 750 1201 774 1232
rect 825 1201 842 1232
rect 900 1201 910 1232
rect 974 1201 978 1232
rect 672 1198 706 1201
rect 740 1198 774 1201
rect 808 1198 842 1201
rect 876 1198 910 1201
rect 944 1198 978 1201
rect 1012 1201 1014 1232
rect 1080 1201 1088 1232
rect 1148 1201 1162 1232
rect 1216 1201 1236 1232
rect 1284 1201 1310 1232
rect 1352 1201 1384 1232
rect 1012 1198 1046 1201
rect 1080 1198 1114 1201
rect 1148 1198 1182 1201
rect 1216 1198 1250 1201
rect 1284 1198 1318 1201
rect 1352 1198 1386 1201
rect 1420 1198 1454 1232
rect 1492 1201 1504 1232
rect 1488 1198 1504 1201
rect 1630 1206 1672 1240
rect 1706 1206 1748 1240
rect 1630 1198 1748 1206
rect 476 1175 510 1196
rect 476 1102 510 1126
rect 1630 1164 1636 1198
rect 1670 1172 1708 1198
rect 1670 1164 1672 1172
rect 1630 1138 1672 1164
rect 1706 1164 1708 1172
rect 1742 1164 1748 1198
rect 1706 1138 1748 1164
rect 1630 1122 1748 1138
rect 1630 1088 1636 1122
rect 1670 1104 1708 1122
rect 1670 1088 1672 1104
rect 476 1029 510 1056
rect 554 1042 570 1076
rect 604 1042 638 1076
rect 672 1042 706 1076
rect 740 1042 774 1076
rect 808 1042 842 1076
rect 876 1042 910 1076
rect 944 1042 978 1076
rect 1012 1042 1046 1076
rect 1080 1042 1114 1076
rect 1158 1042 1182 1076
rect 1236 1042 1250 1076
rect 1314 1042 1318 1076
rect 1352 1042 1358 1076
rect 1420 1042 1435 1076
rect 1488 1042 1512 1076
rect 1630 1070 1672 1088
rect 1706 1088 1708 1104
rect 1742 1088 1748 1122
rect 1706 1070 1748 1088
rect 1630 1046 1748 1070
rect 476 956 510 986
rect 1630 1012 1636 1046
rect 1670 1036 1708 1046
rect 1670 1012 1672 1036
rect 1630 1002 1672 1012
rect 1706 1012 1708 1036
rect 1742 1012 1748 1046
rect 1706 1002 1748 1012
rect 1630 970 1748 1002
rect 1630 936 1636 970
rect 1670 968 1708 970
rect 1670 936 1672 968
rect 1630 934 1672 936
rect 1706 936 1708 968
rect 1742 936 1748 970
rect 1706 934 1748 936
rect 600 920 641 921
rect 675 920 716 921
rect 750 920 791 921
rect 825 920 866 921
rect 900 920 940 921
rect 974 920 1014 921
rect 1048 920 1088 921
rect 1122 920 1162 921
rect 1196 920 1236 921
rect 1270 920 1310 921
rect 1344 920 1384 921
rect 1418 920 1458 921
rect 476 883 510 916
rect 554 887 566 920
rect 554 886 570 887
rect 604 886 638 920
rect 675 887 706 920
rect 750 887 774 920
rect 825 887 842 920
rect 900 887 910 920
rect 974 887 978 920
rect 672 886 706 887
rect 740 886 774 887
rect 808 886 842 887
rect 876 886 910 887
rect 944 886 978 887
rect 1012 887 1014 920
rect 1080 887 1088 920
rect 1148 887 1162 920
rect 1216 887 1236 920
rect 1284 887 1310 920
rect 1352 887 1384 920
rect 1012 886 1046 887
rect 1080 886 1114 887
rect 1148 886 1182 887
rect 1216 886 1250 887
rect 1284 886 1318 887
rect 1352 886 1386 887
rect 1420 886 1454 920
rect 1492 887 1504 920
rect 1488 886 1504 887
rect 1630 900 1748 934
rect 1630 894 1672 900
rect 476 810 510 846
rect 1630 860 1636 894
rect 1670 866 1672 894
rect 1706 894 1748 900
rect 1706 866 1708 894
rect 1670 860 1708 866
rect 1742 860 1748 894
rect 1630 832 1748 860
rect 1630 818 1672 832
rect 476 740 510 776
rect 554 756 566 790
rect 604 756 638 790
rect 675 756 706 790
rect 750 756 774 790
rect 825 756 842 790
rect 900 756 910 790
rect 974 756 978 790
rect 1012 756 1014 790
rect 1080 756 1088 790
rect 1148 756 1162 790
rect 1216 756 1236 790
rect 1284 756 1310 790
rect 1352 756 1384 790
rect 1420 756 1454 790
rect 1492 756 1504 790
rect 1630 784 1636 818
rect 1670 798 1672 818
rect 1706 818 1748 832
rect 1706 798 1708 818
rect 1670 784 1708 798
rect 1742 784 1748 818
rect 1630 764 1748 784
rect 476 669 510 704
rect 1630 741 1672 764
rect 1630 707 1636 741
rect 1670 730 1672 741
rect 1706 741 1748 764
rect 1706 730 1708 741
rect 1670 707 1708 730
rect 1742 707 1748 741
rect 1630 696 1748 707
rect 1630 664 1672 696
rect 476 598 510 632
rect 554 600 570 634
rect 604 600 638 634
rect 672 600 706 634
rect 740 600 774 634
rect 808 600 842 634
rect 876 600 910 634
rect 944 600 978 634
rect 1012 600 1046 634
rect 1080 600 1114 634
rect 1157 600 1182 634
rect 1235 600 1250 634
rect 1313 600 1318 634
rect 1352 600 1357 634
rect 1420 600 1435 634
rect 1488 600 1512 634
rect 1630 630 1636 664
rect 1670 662 1672 664
rect 1706 664 1748 696
rect 1706 662 1708 664
rect 1670 630 1708 662
rect 1742 630 1748 664
rect 1630 628 1748 630
rect 476 522 510 560
rect 1630 594 1672 628
rect 1706 594 1748 628
rect 1630 587 1748 594
rect 1630 553 1636 587
rect 1670 560 1708 587
rect 1670 553 1672 560
rect 1630 526 1672 553
rect 1706 553 1708 560
rect 1742 553 1748 587
rect 1706 526 1748 553
rect 1630 510 1748 526
rect 318 470 436 478
rect 318 436 360 470
rect 394 436 436 470
rect 554 444 566 478
rect 604 444 638 478
rect 675 444 706 478
rect 750 444 774 478
rect 825 444 842 478
rect 900 444 910 478
rect 974 444 978 478
rect 1012 444 1014 478
rect 1080 444 1088 478
rect 1148 444 1162 478
rect 1216 444 1236 478
rect 1284 444 1310 478
rect 1352 444 1384 478
rect 1420 444 1454 478
rect 1492 444 1504 478
rect 1630 476 1636 510
rect 1670 492 1708 510
rect 1670 476 1672 492
rect 1630 458 1672 476
rect 1706 476 1708 492
rect 1742 476 1748 510
rect 1706 458 1748 476
rect 318 402 324 436
rect 358 402 396 436
rect 430 402 436 436
rect 318 362 436 402
rect 1630 433 1748 458
rect 1630 399 1636 433
rect 1670 424 1708 433
rect 1670 399 1672 424
rect 1630 390 1672 399
rect 1706 399 1708 424
rect 1742 399 1748 433
rect 1706 390 1748 399
rect 1630 362 1748 390
rect 318 360 1748 362
rect 318 326 324 360
rect 358 359 1748 360
rect 358 356 425 359
rect 459 356 493 359
rect 527 356 561 359
rect 595 356 629 359
rect 663 356 697 359
rect 731 356 765 359
rect 358 326 396 356
rect 318 322 396 326
rect 459 325 469 356
rect 527 325 542 356
rect 595 325 615 356
rect 663 325 688 356
rect 731 325 761 356
rect 799 325 833 359
rect 867 356 901 359
rect 935 356 969 359
rect 1003 356 1037 359
rect 1071 356 1105 359
rect 1139 356 1173 359
rect 1207 356 1241 359
rect 1275 356 1309 359
rect 868 325 901 356
rect 941 325 969 356
rect 1014 325 1037 356
rect 1087 325 1105 356
rect 1160 325 1173 356
rect 1233 325 1241 356
rect 1306 325 1309 356
rect 1343 356 1377 359
rect 1411 356 1445 359
rect 1479 356 1513 359
rect 1547 356 1581 359
rect 1615 356 1748 359
rect 1343 325 1345 356
rect 1411 325 1418 356
rect 1479 325 1491 356
rect 1547 325 1564 356
rect 430 322 469 325
rect 503 322 542 325
rect 576 322 615 325
rect 649 322 688 325
rect 722 322 761 325
rect 795 322 834 325
rect 868 322 907 325
rect 941 322 980 325
rect 1014 322 1053 325
rect 1087 322 1126 325
rect 1160 322 1199 325
rect 1233 322 1272 325
rect 1306 322 1345 325
rect 1379 322 1418 325
rect 1452 322 1491 325
rect 1525 322 1564 325
rect 318 284 1564 322
rect 318 250 396 284
rect 430 250 469 284
rect 503 250 542 284
rect 576 250 615 284
rect 649 250 688 284
rect 722 250 761 284
rect 795 250 834 284
rect 868 250 907 284
rect 941 250 980 284
rect 1014 250 1053 284
rect 1087 250 1126 284
rect 1160 250 1199 284
rect 1233 250 1272 284
rect 1306 250 1345 284
rect 1379 250 1418 284
rect 1452 250 1491 284
rect 1525 250 1564 284
rect 1670 322 1708 356
rect 1742 322 1748 356
rect 1670 250 1748 322
rect 318 244 1748 250
rect 1898 1400 1904 1434
rect 2010 1400 2016 1434
rect 1898 1359 1906 1400
rect 2008 1359 2016 1400
rect 1898 1325 1904 1359
rect 2010 1325 2016 1359
rect 1898 1284 1906 1325
rect 2008 1284 2016 1325
rect 1898 1250 1904 1284
rect 2010 1250 2016 1284
rect 1898 1209 1906 1250
rect 2008 1209 2016 1250
rect 1898 1175 1904 1209
rect 2010 1175 2016 1209
rect 1898 1134 1906 1175
rect 2008 1134 2016 1175
rect 1898 1100 1904 1134
rect 2010 1100 2016 1134
rect 1898 1059 1906 1100
rect 2008 1059 2016 1100
rect 1898 1025 1904 1059
rect 2010 1025 2016 1059
rect 1898 984 1906 1025
rect 2008 984 2016 1025
rect 1898 950 1904 984
rect 2010 950 2016 984
rect 1898 909 1906 950
rect 2008 909 2016 950
rect 1898 875 1904 909
rect 2010 875 2016 909
rect 1898 835 1906 875
rect 2008 835 2016 875
rect 1898 801 1904 835
rect 2010 801 2016 835
rect 1898 761 1906 801
rect 2008 761 2016 801
rect 1898 727 1904 761
rect 2010 727 2016 761
rect 1898 687 1906 727
rect 2008 687 2016 727
rect 1898 653 1904 687
rect 2010 653 2016 687
rect 1898 613 1906 653
rect 2008 613 2016 653
rect 1898 579 1904 613
rect 2010 579 2016 613
rect 1898 539 1906 579
rect 2008 539 2016 579
rect 1898 505 1904 539
rect 2010 505 2016 539
rect 1898 465 1906 505
rect 2008 465 2016 505
rect 1898 431 1904 465
rect 2010 431 2016 465
rect 1898 391 1906 431
rect 2008 391 2016 431
rect 1898 357 1904 391
rect 2010 357 2016 391
rect 1898 317 1906 357
rect 2008 317 2016 357
rect 1898 283 1904 317
rect 2010 283 2016 317
rect 1898 243 1906 283
rect 2008 243 2016 283
rect 2153 1450 6739 1456
rect 2153 1416 2237 1450
rect 2271 1416 2315 1450
rect 2349 1416 2393 1450
rect 2427 1416 2471 1450
rect 2505 1416 2549 1450
rect 2583 1416 2627 1450
rect 2661 1416 2705 1450
rect 2739 1416 2784 1450
rect 2818 1416 2894 1450
rect 2928 1416 2967 1450
rect 3001 1416 3040 1450
rect 3074 1416 3113 1450
rect 3147 1416 3186 1450
rect 3220 1416 3259 1450
rect 3293 1416 3332 1450
rect 3366 1416 3405 1450
rect 3439 1416 3478 1450
rect 3512 1416 3551 1450
rect 3585 1416 3624 1450
rect 3658 1416 3697 1450
rect 3731 1416 3770 1450
rect 3804 1416 3843 1450
rect 3877 1416 3916 1450
rect 3950 1416 3989 1450
rect 4023 1416 4062 1450
rect 4096 1416 4135 1450
rect 4169 1416 4208 1450
rect 4242 1416 4281 1450
rect 4315 1416 4354 1450
rect 4388 1416 4427 1450
rect 4461 1416 4500 1450
rect 4534 1416 4573 1450
rect 4607 1416 4646 1450
rect 4680 1416 4719 1450
rect 4753 1416 4792 1450
rect 4826 1416 4865 1450
rect 4899 1416 4938 1450
rect 4972 1416 5011 1450
rect 5045 1416 5084 1450
rect 5118 1416 5157 1450
rect 5191 1416 5230 1450
rect 5264 1416 5303 1450
rect 5337 1416 5376 1450
rect 5410 1416 5449 1450
rect 5483 1416 5522 1450
rect 5556 1416 5595 1450
rect 5629 1416 5668 1450
rect 5702 1416 5741 1450
rect 5775 1416 5814 1450
rect 5848 1416 5887 1450
rect 5921 1416 5961 1450
rect 5995 1416 6035 1450
rect 6069 1416 6109 1450
rect 6143 1416 6183 1450
rect 6217 1416 6257 1450
rect 6291 1416 6331 1450
rect 6365 1416 6405 1450
rect 6439 1416 6479 1450
rect 6513 1416 6553 1450
rect 6587 1416 6627 1450
rect 6661 1416 6739 1450
rect 6884 1450 6986 1534
rect 2153 1378 6739 1416
rect 2153 1344 2159 1378
rect 2193 1344 2231 1378
rect 2265 1377 2315 1378
rect 2349 1377 2393 1378
rect 2427 1377 2471 1378
rect 2505 1377 2549 1378
rect 2583 1377 2627 1378
rect 2661 1377 2705 1378
rect 2739 1377 2784 1378
rect 2818 1377 2894 1378
rect 2928 1377 2967 1378
rect 3001 1377 3040 1378
rect 3074 1377 3113 1378
rect 3147 1377 3186 1378
rect 3220 1377 3259 1378
rect 3293 1377 3332 1378
rect 3366 1377 3405 1378
rect 3439 1377 3478 1378
rect 3512 1377 3551 1378
rect 3585 1377 3624 1378
rect 3658 1377 3697 1378
rect 3731 1377 3770 1378
rect 3804 1377 3843 1378
rect 3877 1377 3916 1378
rect 3950 1377 3989 1378
rect 4023 1377 4062 1378
rect 4096 1377 4135 1378
rect 4169 1377 4208 1378
rect 4242 1377 4281 1378
rect 4315 1377 4354 1378
rect 4388 1377 4427 1378
rect 2265 1344 2287 1377
rect 2349 1344 2355 1377
rect 2153 1343 2287 1344
rect 2321 1343 2355 1344
rect 2389 1344 2393 1377
rect 2457 1344 2471 1377
rect 2525 1344 2549 1377
rect 2389 1343 2423 1344
rect 2457 1343 2491 1344
rect 2525 1343 2559 1344
rect 2593 1343 2627 1377
rect 2661 1343 2695 1377
rect 2739 1344 2763 1377
rect 2818 1344 2831 1377
rect 2729 1343 2763 1344
rect 2797 1343 2831 1344
rect 2865 1344 2894 1377
rect 2865 1343 2899 1344
rect 2933 1343 2967 1377
rect 3001 1343 3035 1377
rect 3074 1344 3103 1377
rect 3147 1344 3171 1377
rect 3220 1344 3239 1377
rect 3293 1344 3307 1377
rect 3366 1344 3375 1377
rect 3439 1344 3443 1377
rect 3069 1343 3103 1344
rect 3137 1343 3171 1344
rect 3205 1343 3239 1344
rect 3273 1343 3307 1344
rect 3341 1343 3375 1344
rect 3409 1343 3443 1344
rect 3477 1344 3478 1377
rect 3545 1344 3551 1377
rect 3613 1344 3624 1377
rect 3681 1344 3697 1377
rect 3749 1344 3770 1377
rect 3817 1344 3843 1377
rect 3885 1344 3916 1377
rect 3477 1343 3511 1344
rect 3545 1343 3579 1344
rect 3613 1343 3647 1344
rect 3681 1343 3715 1344
rect 3749 1343 3783 1344
rect 3817 1343 3851 1344
rect 3885 1343 3919 1344
rect 3953 1343 3987 1377
rect 4023 1344 4055 1377
rect 4096 1344 4123 1377
rect 4169 1344 4191 1377
rect 4242 1344 4259 1377
rect 4315 1344 4327 1377
rect 4388 1344 4395 1377
rect 4461 1344 4500 1378
rect 4534 1377 4573 1378
rect 4607 1377 4646 1378
rect 4680 1377 4719 1378
rect 4753 1377 4792 1378
rect 4826 1377 4865 1378
rect 4899 1377 4938 1378
rect 4972 1377 5011 1378
rect 5045 1377 5084 1378
rect 5118 1377 5157 1378
rect 5191 1377 5230 1378
rect 5264 1377 5303 1378
rect 5337 1377 5376 1378
rect 5410 1377 5449 1378
rect 5483 1377 5522 1378
rect 5556 1377 5595 1378
rect 5629 1377 5668 1378
rect 5702 1377 5741 1378
rect 5775 1377 5814 1378
rect 5848 1377 5887 1378
rect 5921 1377 5961 1378
rect 5995 1377 6035 1378
rect 6069 1377 6109 1378
rect 6143 1377 6183 1378
rect 6217 1377 6257 1378
rect 6291 1377 6331 1378
rect 6365 1377 6405 1378
rect 6439 1377 6479 1378
rect 6513 1377 6553 1378
rect 6587 1377 6627 1378
rect 4534 1344 4558 1377
rect 4607 1344 4626 1377
rect 4680 1344 4694 1377
rect 4753 1344 4762 1377
rect 4826 1344 4830 1377
rect 4021 1343 4055 1344
rect 4089 1343 4123 1344
rect 4157 1343 4191 1344
rect 4225 1343 4259 1344
rect 4293 1343 4327 1344
rect 4361 1343 4395 1344
rect 4429 1343 4558 1344
rect 4592 1343 4626 1344
rect 4660 1343 4694 1344
rect 4728 1343 4762 1344
rect 4796 1343 4830 1344
rect 4864 1344 4865 1377
rect 4932 1344 4938 1377
rect 5000 1344 5011 1377
rect 5068 1344 5084 1377
rect 5136 1344 5157 1377
rect 5204 1344 5230 1377
rect 5272 1344 5303 1377
rect 4864 1343 4898 1344
rect 4932 1343 4966 1344
rect 5000 1343 5034 1344
rect 5068 1343 5102 1344
rect 5136 1343 5170 1344
rect 5204 1343 5238 1344
rect 5272 1343 5306 1344
rect 5340 1343 5374 1377
rect 5410 1344 5442 1377
rect 5483 1344 5510 1377
rect 5556 1344 5578 1377
rect 5629 1344 5646 1377
rect 5702 1344 5714 1377
rect 5775 1344 5782 1377
rect 5848 1344 5850 1377
rect 5408 1343 5442 1344
rect 5476 1343 5510 1344
rect 5544 1343 5578 1344
rect 5612 1343 5646 1344
rect 5680 1343 5714 1344
rect 5748 1343 5782 1344
rect 5816 1343 5850 1344
rect 5884 1344 5887 1377
rect 5952 1344 5961 1377
rect 6020 1344 6035 1377
rect 6088 1344 6109 1377
rect 6156 1344 6183 1377
rect 6224 1344 6257 1377
rect 5884 1343 5918 1344
rect 5952 1343 5986 1344
rect 6020 1343 6054 1344
rect 6088 1343 6122 1344
rect 6156 1343 6190 1344
rect 6224 1343 6258 1344
rect 6292 1343 6326 1377
rect 6365 1344 6394 1377
rect 6439 1344 6462 1377
rect 6513 1344 6530 1377
rect 6587 1344 6598 1377
rect 6360 1343 6394 1344
rect 6428 1343 6462 1344
rect 6496 1343 6530 1344
rect 6564 1343 6598 1344
rect 2153 1338 6627 1343
rect 2153 1312 2271 1338
rect 2153 1305 2195 1312
rect 2153 1271 2159 1305
rect 2193 1278 2195 1305
rect 2229 1305 2271 1312
rect 2229 1278 2231 1305
rect 2193 1271 2231 1278
rect 2265 1271 2271 1305
rect 2153 1244 2271 1271
rect 2153 1232 2195 1244
rect 2153 1198 2159 1232
rect 2193 1210 2195 1232
rect 2229 1232 2271 1244
rect 2229 1210 2231 1232
rect 2193 1198 2231 1210
rect 2265 1198 2271 1232
rect 2389 1224 2401 1258
rect 2439 1224 2473 1258
rect 2509 1224 2541 1258
rect 2583 1224 2609 1258
rect 2657 1224 2677 1258
rect 2731 1224 2745 1258
rect 2805 1224 2813 1258
rect 2879 1224 2881 1258
rect 2915 1224 2919 1258
rect 2983 1224 2993 1258
rect 3051 1224 3067 1258
rect 3119 1224 3141 1258
rect 3187 1224 3215 1258
rect 3255 1224 3289 1258
rect 3323 1224 3357 1258
rect 3397 1224 3425 1258
rect 3471 1224 3493 1258
rect 3544 1224 3561 1258
rect 3617 1224 3629 1258
rect 3690 1224 3697 1258
rect 3763 1224 3765 1258
rect 3799 1224 3802 1258
rect 3867 1224 3875 1258
rect 3935 1224 3948 1258
rect 4003 1224 4021 1258
rect 4071 1224 4094 1258
rect 4139 1224 4167 1258
rect 4207 1224 4240 1258
rect 4275 1224 4309 1258
rect 4347 1224 4359 1258
rect 4533 1224 4545 1258
rect 4583 1224 4617 1258
rect 4652 1224 4685 1258
rect 4725 1224 4753 1258
rect 4798 1224 4821 1258
rect 4871 1224 4889 1258
rect 4944 1224 4957 1258
rect 5017 1224 5025 1258
rect 5090 1224 5093 1258
rect 5127 1224 5129 1258
rect 5195 1224 5202 1258
rect 5263 1224 5275 1258
rect 5331 1224 5348 1258
rect 5399 1224 5421 1258
rect 5467 1224 5495 1258
rect 5535 1224 5569 1258
rect 5603 1224 5637 1258
rect 5677 1224 5705 1258
rect 5751 1224 5773 1258
rect 5825 1224 5841 1258
rect 5899 1224 5909 1258
rect 5973 1224 5977 1258
rect 6011 1224 6013 1258
rect 6079 1224 6087 1258
rect 6147 1224 6161 1258
rect 6215 1224 6235 1258
rect 6283 1224 6309 1258
rect 6351 1224 6383 1258
rect 6419 1224 6453 1258
rect 6491 1224 6503 1258
rect 2153 1176 2271 1198
rect 2153 1159 2195 1176
rect 2153 1125 2159 1159
rect 2193 1142 2195 1159
rect 2229 1159 2271 1176
rect 2229 1142 2231 1159
rect 2193 1125 2231 1142
rect 2265 1125 2271 1159
rect 2153 1108 2271 1125
rect 2153 1086 2195 1108
rect 2153 1052 2159 1086
rect 2193 1074 2195 1086
rect 2229 1086 2271 1108
rect 2229 1074 2231 1086
rect 2193 1052 2231 1074
rect 2265 1052 2271 1086
rect 2153 1040 2271 1052
rect 2153 1013 2195 1040
rect 2153 979 2159 1013
rect 2193 1006 2195 1013
rect 2229 1013 2271 1040
rect 2229 1006 2231 1013
rect 2193 979 2231 1006
rect 2265 979 2271 1013
rect 2153 972 2271 979
rect 2153 940 2195 972
rect 2153 906 2159 940
rect 2193 938 2195 940
rect 2229 940 2271 972
rect 2229 938 2231 940
rect 2193 906 2231 938
rect 2265 906 2271 940
rect 2153 904 2271 906
rect 2153 870 2195 904
rect 2229 870 2271 904
rect 2153 867 2271 870
rect 2153 833 2159 867
rect 2193 836 2231 867
rect 2193 833 2195 836
rect 2153 802 2195 833
rect 2229 833 2231 836
rect 2265 833 2271 867
rect 2229 802 2271 833
rect 2153 794 2271 802
rect 2153 760 2159 794
rect 2193 768 2231 794
rect 2193 760 2195 768
rect 2153 734 2195 760
rect 2229 760 2231 768
rect 2265 760 2271 794
rect 2229 734 2271 760
rect 2153 721 2271 734
rect 2153 687 2159 721
rect 2193 700 2231 721
rect 2193 687 2195 700
rect 2153 666 2195 687
rect 2229 687 2231 700
rect 2265 687 2271 721
rect 2229 666 2271 687
rect 2153 648 2271 666
rect 2153 614 2159 648
rect 2193 632 2231 648
rect 2193 614 2195 632
rect 2153 598 2195 614
rect 2229 614 2231 632
rect 2265 614 2271 648
rect 2229 598 2271 614
rect 2153 575 2271 598
rect 2153 541 2159 575
rect 2193 564 2231 575
rect 2193 541 2195 564
rect 2153 530 2195 541
rect 2229 541 2231 564
rect 2265 541 2271 575
rect 2311 1201 2345 1213
rect 2311 1128 2345 1163
rect 6547 1201 6581 1213
rect 6547 1129 6581 1163
rect 2311 1055 2345 1089
rect 2389 1068 2401 1102
rect 2439 1068 2473 1102
rect 2509 1068 2541 1102
rect 2583 1068 2609 1102
rect 2657 1068 2677 1102
rect 2731 1068 2745 1102
rect 2805 1068 2813 1102
rect 2879 1068 2881 1102
rect 2915 1068 2919 1102
rect 2983 1068 2993 1102
rect 3051 1068 3067 1102
rect 3119 1068 3141 1102
rect 3187 1068 3215 1102
rect 3255 1068 3289 1102
rect 3323 1068 3357 1102
rect 3397 1068 3425 1102
rect 3471 1068 3493 1102
rect 3544 1068 3561 1102
rect 3617 1068 3629 1102
rect 3690 1068 3697 1102
rect 3763 1068 3765 1102
rect 3799 1068 3802 1102
rect 3867 1068 3875 1102
rect 3935 1068 3948 1102
rect 4003 1068 4021 1102
rect 4071 1068 4094 1102
rect 4139 1068 4167 1102
rect 4207 1068 4240 1102
rect 4275 1068 4309 1102
rect 4347 1068 4359 1102
rect 4533 1068 4545 1102
rect 4583 1068 4617 1102
rect 4652 1068 4685 1102
rect 4725 1068 4753 1102
rect 4798 1068 4821 1102
rect 4871 1068 4889 1102
rect 4944 1068 4957 1102
rect 5017 1068 5025 1102
rect 5090 1068 5093 1102
rect 5127 1068 5129 1102
rect 5195 1068 5202 1102
rect 5263 1068 5275 1102
rect 5331 1068 5348 1102
rect 5399 1068 5421 1102
rect 5467 1068 5495 1102
rect 5535 1068 5569 1102
rect 5603 1068 5637 1102
rect 5677 1068 5705 1102
rect 5751 1068 5773 1102
rect 5825 1068 5841 1102
rect 5899 1068 5909 1102
rect 5973 1068 5977 1102
rect 6011 1068 6013 1102
rect 6079 1068 6087 1102
rect 6147 1068 6161 1102
rect 6215 1068 6235 1102
rect 6283 1068 6309 1102
rect 6351 1068 6383 1102
rect 6419 1068 6453 1102
rect 6491 1068 6503 1102
rect 2311 981 2345 1015
rect 6547 1056 6581 1089
rect 6547 983 6581 1015
rect 2311 907 2345 940
rect 2389 912 2401 946
rect 2439 912 2473 946
rect 2509 912 2541 946
rect 2583 912 2609 946
rect 2657 912 2677 946
rect 2731 912 2745 946
rect 2805 912 2813 946
rect 2879 912 2881 946
rect 2915 912 2919 946
rect 2983 912 2993 946
rect 3051 912 3067 946
rect 3119 912 3141 946
rect 3187 912 3215 946
rect 3255 912 3289 946
rect 3323 912 3357 946
rect 3397 912 3425 946
rect 3471 912 3493 946
rect 3544 912 3561 946
rect 3617 912 3629 946
rect 3690 912 3697 946
rect 3763 912 3765 946
rect 3799 912 3802 946
rect 3867 912 3875 946
rect 3935 912 3948 946
rect 4003 912 4021 946
rect 4071 912 4094 946
rect 4139 912 4167 946
rect 4207 912 4240 946
rect 4275 912 4309 946
rect 4347 912 4359 946
rect 4533 912 4545 946
rect 4583 912 4617 946
rect 4652 912 4685 946
rect 4725 912 4753 946
rect 4798 912 4821 946
rect 4871 912 4889 946
rect 4944 912 4957 946
rect 5017 912 5025 946
rect 5090 912 5093 946
rect 5127 912 5129 946
rect 5195 912 5202 946
rect 5263 912 5275 946
rect 5331 912 5348 946
rect 5399 912 5421 946
rect 5467 912 5495 946
rect 5535 912 5569 946
rect 5603 912 5637 946
rect 5677 912 5705 946
rect 5751 912 5773 946
rect 5825 912 5841 946
rect 5899 912 5909 946
rect 5973 912 5977 946
rect 6011 912 6013 946
rect 6079 912 6087 946
rect 6147 912 6161 946
rect 6215 912 6235 946
rect 6283 912 6309 946
rect 6351 912 6383 946
rect 6419 912 6453 946
rect 6491 912 6503 946
rect 2311 833 2345 865
rect 6547 910 6581 940
rect 6547 837 6581 865
rect 2311 759 2345 790
rect 2389 756 2401 790
rect 2439 756 2473 790
rect 2509 756 2541 790
rect 2583 756 2609 790
rect 2657 756 2677 790
rect 2731 756 2745 790
rect 2805 756 2813 790
rect 2879 756 2881 790
rect 2915 756 2919 790
rect 2983 756 2993 790
rect 3051 756 3067 790
rect 3119 756 3141 790
rect 3187 756 3215 790
rect 3255 756 3289 790
rect 3323 756 3357 790
rect 3397 756 3425 790
rect 3471 756 3493 790
rect 3544 756 3561 790
rect 3617 756 3629 790
rect 3690 756 3697 790
rect 3763 756 3765 790
rect 3799 756 3802 790
rect 3867 756 3875 790
rect 3935 756 3948 790
rect 4003 756 4021 790
rect 4071 756 4094 790
rect 4139 756 4167 790
rect 4207 756 4240 790
rect 4275 756 4309 790
rect 4347 756 4359 790
rect 4533 756 4545 790
rect 4583 756 4617 790
rect 4652 756 4685 790
rect 4725 756 4753 790
rect 4798 756 4821 790
rect 4871 756 4889 790
rect 4944 756 4957 790
rect 5017 756 5025 790
rect 5090 756 5093 790
rect 5127 756 5129 790
rect 5195 756 5202 790
rect 5263 756 5275 790
rect 5331 756 5348 790
rect 5399 756 5421 790
rect 5467 756 5495 790
rect 5535 756 5569 790
rect 5603 756 5637 790
rect 5677 756 5705 790
rect 5751 756 5773 790
rect 5825 756 5841 790
rect 5899 756 5909 790
rect 5973 756 5977 790
rect 6011 756 6013 790
rect 6079 756 6087 790
rect 6147 756 6161 790
rect 6215 756 6235 790
rect 6283 756 6309 790
rect 6351 756 6383 790
rect 6419 756 6453 790
rect 6491 756 6503 790
rect 6547 764 6581 790
rect 2311 685 2345 715
rect 2311 599 2345 640
rect 6547 691 6581 715
rect 2389 600 2401 634
rect 2439 600 2473 634
rect 2509 600 2541 634
rect 2583 600 2609 634
rect 2657 600 2677 634
rect 2731 600 2745 634
rect 2805 600 2813 634
rect 2879 600 2881 634
rect 2915 600 2919 634
rect 2983 600 2993 634
rect 3051 600 3067 634
rect 3119 600 3141 634
rect 3187 600 3215 634
rect 3255 600 3289 634
rect 3323 600 3357 634
rect 3397 600 3425 634
rect 3471 600 3493 634
rect 3544 600 3561 634
rect 3617 600 3629 634
rect 3690 600 3697 634
rect 3763 600 3765 634
rect 3799 600 3802 634
rect 3867 600 3875 634
rect 3935 600 3948 634
rect 4003 600 4021 634
rect 4071 600 4094 634
rect 4139 600 4167 634
rect 4207 600 4240 634
rect 4275 600 4309 634
rect 4347 600 4359 634
rect 4533 600 4545 634
rect 4583 600 4617 634
rect 4652 600 4685 634
rect 4725 600 4753 634
rect 4798 600 4821 634
rect 4871 600 4889 634
rect 4944 600 4957 634
rect 5017 600 5025 634
rect 5090 600 5093 634
rect 5127 600 5129 634
rect 5195 600 5202 634
rect 5263 600 5275 634
rect 5331 600 5348 634
rect 5399 600 5421 634
rect 5467 600 5495 634
rect 5535 600 5569 634
rect 5603 600 5637 634
rect 5677 600 5705 634
rect 5751 600 5773 634
rect 5825 600 5841 634
rect 5899 600 5909 634
rect 5973 600 5977 634
rect 6011 600 6013 634
rect 6079 600 6087 634
rect 6147 600 6161 634
rect 6215 600 6235 634
rect 6283 600 6309 634
rect 6351 600 6383 634
rect 6419 600 6453 634
rect 6491 600 6503 634
rect 2311 549 2345 565
rect 6547 599 6581 640
rect 6547 549 6581 565
rect 6621 1200 6627 1338
rect 6733 1200 6739 1378
rect 6621 1172 6739 1200
rect 6621 1161 6663 1172
rect 6621 1127 6627 1161
rect 6661 1138 6663 1161
rect 6697 1161 6739 1172
rect 6697 1138 6699 1161
rect 6661 1127 6699 1138
rect 6733 1127 6739 1161
rect 6621 1104 6739 1127
rect 6621 1088 6663 1104
rect 6621 1054 6627 1088
rect 6661 1070 6663 1088
rect 6697 1088 6739 1104
rect 6697 1070 6699 1088
rect 6661 1054 6699 1070
rect 6733 1054 6739 1088
rect 6621 1036 6739 1054
rect 6621 1015 6663 1036
rect 6621 981 6627 1015
rect 6661 1002 6663 1015
rect 6697 1015 6739 1036
rect 6697 1002 6699 1015
rect 6661 981 6699 1002
rect 6733 981 6739 1015
rect 6621 968 6739 981
rect 6621 942 6663 968
rect 6621 908 6627 942
rect 6661 934 6663 942
rect 6697 942 6739 968
rect 6697 934 6699 942
rect 6661 908 6699 934
rect 6733 908 6739 942
rect 6621 900 6739 908
rect 6621 869 6663 900
rect 6621 835 6627 869
rect 6661 866 6663 869
rect 6697 869 6739 900
rect 6697 866 6699 869
rect 6661 835 6699 866
rect 6733 835 6739 869
rect 6621 832 6739 835
rect 6621 798 6663 832
rect 6697 798 6739 832
rect 6621 796 6739 798
rect 6621 762 6627 796
rect 6661 764 6699 796
rect 6661 762 6663 764
rect 6621 730 6663 762
rect 6697 762 6699 764
rect 6733 762 6739 796
rect 6697 730 6739 762
rect 6621 723 6739 730
rect 6621 689 6627 723
rect 6661 696 6699 723
rect 6661 689 6663 696
rect 6621 662 6663 689
rect 6697 689 6699 696
rect 6733 689 6739 723
rect 6697 662 6739 689
rect 6621 650 6739 662
rect 6621 616 6627 650
rect 6661 628 6699 650
rect 6661 616 6663 628
rect 6621 594 6663 616
rect 6697 616 6699 628
rect 6733 616 6739 650
rect 6697 594 6739 616
rect 6621 577 6739 594
rect 2229 530 2271 541
rect 2153 502 2271 530
rect 2153 324 2159 502
rect 2265 364 2271 502
rect 6621 543 6627 577
rect 6661 560 6699 577
rect 6661 543 6663 560
rect 6621 526 6663 543
rect 6697 543 6699 560
rect 6733 543 6739 577
rect 6697 526 6739 543
rect 6621 504 6739 526
rect 2389 444 2401 478
rect 2439 444 2473 478
rect 2509 444 2541 478
rect 2583 444 2609 478
rect 2657 444 2677 478
rect 2731 444 2745 478
rect 2805 444 2813 478
rect 2879 444 2881 478
rect 2915 444 2919 478
rect 2983 444 2993 478
rect 3051 444 3067 478
rect 3119 444 3141 478
rect 3187 444 3215 478
rect 3255 444 3289 478
rect 3323 444 3357 478
rect 3397 444 3425 478
rect 3471 444 3493 478
rect 3544 444 3561 478
rect 3617 444 3629 478
rect 3690 444 3697 478
rect 3763 444 3765 478
rect 3799 444 3802 478
rect 3867 444 3875 478
rect 3935 444 3948 478
rect 4003 444 4021 478
rect 4071 444 4094 478
rect 4139 444 4167 478
rect 4207 444 4240 478
rect 4275 444 4309 478
rect 4347 444 4359 478
rect 4533 444 4545 478
rect 4583 444 4617 478
rect 4652 444 4685 478
rect 4725 444 4753 478
rect 4798 444 4821 478
rect 4871 444 4889 478
rect 4944 444 4957 478
rect 5017 444 5025 478
rect 5090 444 5093 478
rect 5127 444 5129 478
rect 5195 444 5202 478
rect 5263 444 5275 478
rect 5331 444 5348 478
rect 5399 444 5421 478
rect 5467 444 5495 478
rect 5535 444 5569 478
rect 5603 444 5637 478
rect 5677 444 5705 478
rect 5751 444 5773 478
rect 5825 444 5841 478
rect 5899 444 5909 478
rect 5973 444 5977 478
rect 6011 444 6013 478
rect 6079 444 6087 478
rect 6147 444 6161 478
rect 6215 444 6235 478
rect 6283 444 6309 478
rect 6351 444 6383 478
rect 6419 444 6453 478
rect 6491 444 6503 478
rect 6621 470 6627 504
rect 6661 492 6699 504
rect 6661 470 6663 492
rect 6621 458 6663 470
rect 6697 470 6699 492
rect 6733 470 6739 504
rect 6697 458 6739 470
rect 6621 431 6739 458
rect 6621 397 6627 431
rect 6661 424 6699 431
rect 6661 397 6663 424
rect 6621 390 6663 397
rect 6697 397 6699 424
rect 6733 397 6739 431
rect 6697 390 6739 397
rect 6621 364 6739 390
rect 2265 359 6739 364
rect 2294 358 2328 359
rect 2362 358 2396 359
rect 2430 358 2464 359
rect 2498 358 2532 359
rect 2566 358 2600 359
rect 2634 358 2668 359
rect 2702 358 2736 359
rect 2770 358 2804 359
rect 2838 358 2872 359
rect 2906 358 2940 359
rect 2974 358 3008 359
rect 3042 358 3076 359
rect 3110 358 3144 359
rect 3178 358 3212 359
rect 3246 358 3280 359
rect 3314 358 3348 359
rect 3382 358 3416 359
rect 3450 358 3484 359
rect 3518 358 3552 359
rect 3586 358 3620 359
rect 3654 358 3688 359
rect 3722 358 3756 359
rect 3790 358 3824 359
rect 3858 358 3892 359
rect 3926 358 3960 359
rect 3994 358 4028 359
rect 4062 358 4096 359
rect 4130 358 4164 359
rect 4198 358 4232 359
rect 4266 358 4300 359
rect 4334 358 4368 359
rect 4402 358 4436 359
rect 4470 358 4504 359
rect 4538 358 4572 359
rect 4606 358 4640 359
rect 4674 358 4708 359
rect 4742 358 4776 359
rect 4810 358 4844 359
rect 4878 358 4912 359
rect 4946 358 4980 359
rect 5014 358 5048 359
rect 5082 358 5116 359
rect 5150 358 5184 359
rect 5218 358 5252 359
rect 5286 358 5320 359
rect 5354 358 5388 359
rect 5422 358 5456 359
rect 5490 358 5524 359
rect 5558 358 5592 359
rect 5626 358 5660 359
rect 5694 358 5728 359
rect 5762 358 5796 359
rect 5830 358 5864 359
rect 5898 358 5932 359
rect 5966 358 6000 359
rect 6034 358 6068 359
rect 6102 358 6136 359
rect 6170 358 6204 359
rect 6238 358 6272 359
rect 6306 358 6340 359
rect 6374 358 6408 359
rect 6442 358 6476 359
rect 6510 358 6544 359
rect 6578 358 6739 359
rect 2294 325 2304 358
rect 2362 325 2377 358
rect 2430 325 2450 358
rect 2498 325 2523 358
rect 2265 324 2304 325
rect 2338 324 2377 325
rect 2411 324 2450 325
rect 2484 324 2523 325
rect 2153 286 2523 324
rect 2153 252 2231 286
rect 2265 252 2304 286
rect 2338 252 2377 286
rect 2411 252 2450 286
rect 2484 252 2523 286
rect 6661 324 6699 358
rect 6733 324 6739 358
rect 6661 252 6739 324
rect 2153 246 6739 252
rect 6876 1416 6884 1448
rect 7157 1450 11757 1456
rect 6986 1416 6994 1448
rect 6876 1382 6882 1416
rect 6988 1382 6994 1416
rect 6876 1343 6884 1382
rect 6986 1343 6994 1382
rect 6876 1309 6882 1343
rect 6988 1309 6994 1343
rect 6876 1270 6884 1309
rect 6986 1270 6994 1309
rect 6876 1236 6882 1270
rect 6988 1236 6994 1270
rect 6876 1197 6884 1236
rect 6986 1197 6994 1236
rect 6876 1163 6882 1197
rect 6988 1163 6994 1197
rect 6876 1124 6884 1163
rect 6986 1124 6994 1163
rect 6876 1090 6882 1124
rect 6988 1090 6994 1124
rect 6876 1051 6884 1090
rect 6986 1051 6994 1090
rect 6876 1017 6882 1051
rect 6988 1017 6994 1051
rect 6876 978 6884 1017
rect 6986 978 6994 1017
rect 6876 944 6882 978
rect 6988 944 6994 978
rect 6876 905 6884 944
rect 6986 905 6994 944
rect 6876 871 6882 905
rect 6988 871 6994 905
rect 6876 832 6884 871
rect 6986 832 6994 871
rect 6876 798 6882 832
rect 6988 798 6994 832
rect 6876 759 6884 798
rect 6986 759 6994 798
rect 6876 725 6882 759
rect 6988 725 6994 759
rect 6876 686 6884 725
rect 6986 686 6994 725
rect 6876 652 6882 686
rect 6988 652 6994 686
rect 6876 613 6884 652
rect 6986 613 6994 652
rect 6876 579 6882 613
rect 6988 579 6994 613
rect 6876 539 6884 579
rect 6986 539 6994 579
rect 6876 505 6882 539
rect 6988 505 6994 539
rect 6876 465 6884 505
rect 6986 465 6994 505
rect 6876 431 6882 465
rect 6988 431 6994 465
rect 6876 391 6884 431
rect 6986 391 6994 431
rect 6876 357 6882 391
rect 6988 357 6994 391
rect 6876 317 6884 357
rect 6986 317 6994 357
rect 6876 283 6882 317
rect 6988 283 6994 317
rect 6876 260 6884 283
rect 6986 260 6994 283
rect 1898 209 1904 243
rect 2010 209 2016 243
rect 1898 177 1906 209
rect 167 171 1906 177
rect 2008 177 2016 209
rect 6876 243 6994 260
rect 7157 1416 7241 1450
rect 7275 1416 7319 1450
rect 7353 1416 7397 1450
rect 7431 1416 7475 1450
rect 7509 1416 7553 1450
rect 7587 1416 7631 1450
rect 7665 1416 7709 1450
rect 7743 1416 7788 1450
rect 7822 1416 7898 1450
rect 7157 1378 7898 1416
rect 7157 1344 7163 1378
rect 7197 1344 7235 1378
rect 7269 1377 7319 1378
rect 7353 1377 7397 1378
rect 7431 1377 7475 1378
rect 7509 1377 7553 1378
rect 7587 1377 7631 1378
rect 7665 1377 7709 1378
rect 7743 1377 7788 1378
rect 7822 1377 7898 1378
rect 11460 1416 11499 1450
rect 11533 1416 11572 1450
rect 11606 1416 11645 1450
rect 11679 1416 11757 1450
rect 11460 1378 11757 1416
rect 11460 1377 11499 1378
rect 11533 1377 11572 1378
rect 11606 1377 11645 1378
rect 7298 1344 7319 1377
rect 7366 1344 7397 1377
rect 7157 1343 7264 1344
rect 7298 1343 7332 1344
rect 7366 1343 7400 1344
rect 7434 1343 7468 1377
rect 7509 1344 7536 1377
rect 7587 1344 7604 1377
rect 7665 1344 7672 1377
rect 7502 1343 7536 1344
rect 7570 1343 7604 1344
rect 7638 1343 7672 1344
rect 7706 1344 7709 1377
rect 7774 1344 7788 1377
rect 7706 1343 7740 1344
rect 7774 1343 7808 1344
rect 7842 1343 7876 1377
rect 11460 1344 11472 1377
rect 11533 1344 11540 1377
rect 11606 1344 11608 1377
rect 7910 1343 7944 1344
rect 7978 1343 8012 1344
rect 8046 1343 8080 1344
rect 8114 1343 8148 1344
rect 8182 1343 8216 1344
rect 8250 1343 8284 1344
rect 8318 1343 8352 1344
rect 8386 1343 8420 1344
rect 8454 1343 8488 1344
rect 8522 1343 8556 1344
rect 8590 1343 8624 1344
rect 8658 1343 8692 1344
rect 8726 1343 8760 1344
rect 8794 1343 8828 1344
rect 8862 1343 8896 1344
rect 8930 1343 8964 1344
rect 8998 1343 9032 1344
rect 9066 1343 9100 1344
rect 9134 1343 9168 1344
rect 9202 1343 9236 1344
rect 9270 1343 9304 1344
rect 9338 1343 9372 1344
rect 9406 1343 9500 1344
rect 9534 1343 9568 1344
rect 9602 1343 9636 1344
rect 9670 1343 9704 1344
rect 9738 1343 9772 1344
rect 9806 1343 9840 1344
rect 9874 1343 9908 1344
rect 9942 1343 9976 1344
rect 10010 1343 10044 1344
rect 10078 1343 10112 1344
rect 10146 1343 10180 1344
rect 10214 1343 10248 1344
rect 10282 1343 10316 1344
rect 10350 1343 10384 1344
rect 10418 1343 10452 1344
rect 10486 1343 10520 1344
rect 10554 1343 10588 1344
rect 10622 1343 10656 1344
rect 10690 1343 10724 1344
rect 10758 1343 10792 1344
rect 10826 1343 10860 1344
rect 10894 1343 10928 1344
rect 10962 1343 10996 1344
rect 11030 1343 11064 1344
rect 11098 1343 11132 1344
rect 11166 1343 11200 1344
rect 11234 1343 11268 1344
rect 11302 1343 11336 1344
rect 11370 1343 11404 1344
rect 11438 1343 11472 1344
rect 11506 1343 11540 1344
rect 11574 1343 11608 1344
rect 11642 1343 11645 1377
rect 7157 1338 11645 1343
rect 7157 1308 7275 1338
rect 7157 1305 7199 1308
rect 7157 1271 7163 1305
rect 7197 1274 7199 1305
rect 7233 1305 7275 1308
rect 7233 1274 7235 1305
rect 7197 1271 7235 1274
rect 7269 1271 7275 1305
rect 7157 1240 7275 1271
rect 7157 1232 7199 1240
rect 7157 1198 7163 1232
rect 7197 1206 7199 1232
rect 7233 1232 7275 1240
rect 7233 1206 7235 1232
rect 7197 1198 7235 1206
rect 7269 1198 7275 1232
rect 7454 1224 7462 1258
rect 7528 1224 7530 1258
rect 7564 1224 7568 1258
rect 7632 1224 7642 1258
rect 7700 1224 7716 1258
rect 7768 1224 7790 1258
rect 7836 1224 7864 1258
rect 7904 1224 7938 1258
rect 7972 1224 8006 1258
rect 8046 1224 8074 1258
rect 8120 1224 8142 1258
rect 8194 1224 8210 1258
rect 8268 1224 8278 1258
rect 8342 1224 8346 1258
rect 8380 1224 8382 1258
rect 8448 1224 8456 1258
rect 8516 1224 8529 1258
rect 8584 1224 8602 1258
rect 8652 1224 8675 1258
rect 8720 1224 8748 1258
rect 8788 1224 8821 1258
rect 8856 1224 8890 1258
rect 8928 1224 8958 1258
rect 9001 1224 9026 1258
rect 9074 1224 9094 1258
rect 9147 1224 9162 1258
rect 9220 1224 9230 1258
rect 9293 1224 9298 1258
rect 9400 1224 9416 1258
rect 9552 1224 9564 1258
rect 9602 1224 9636 1258
rect 9671 1224 9704 1258
rect 9744 1224 9772 1258
rect 9817 1224 9840 1258
rect 9890 1224 9908 1258
rect 9963 1224 9976 1258
rect 10036 1224 10044 1258
rect 10109 1224 10112 1258
rect 10146 1224 10148 1258
rect 10214 1224 10221 1258
rect 10282 1224 10294 1258
rect 10350 1224 10367 1258
rect 10418 1224 10440 1258
rect 10486 1224 10514 1258
rect 10554 1224 10588 1258
rect 10622 1224 10656 1258
rect 10696 1224 10724 1258
rect 10770 1224 10792 1258
rect 10844 1224 10860 1258
rect 10918 1224 10928 1258
rect 10992 1224 10996 1258
rect 11030 1224 11032 1258
rect 11098 1224 11106 1258
rect 11166 1224 11180 1258
rect 11234 1224 11254 1258
rect 11302 1224 11328 1258
rect 11370 1224 11402 1258
rect 11438 1224 11472 1258
rect 11510 1224 11522 1258
rect 7157 1172 7275 1198
rect 7157 1159 7199 1172
rect 7157 1125 7163 1159
rect 7197 1138 7199 1159
rect 7233 1159 7275 1172
rect 7233 1138 7235 1159
rect 7197 1125 7235 1138
rect 7269 1125 7275 1159
rect 7157 1104 7275 1125
rect 7157 1086 7199 1104
rect 7157 1052 7163 1086
rect 7197 1070 7199 1086
rect 7233 1086 7275 1104
rect 7233 1070 7235 1086
rect 7197 1052 7235 1070
rect 7269 1052 7275 1086
rect 7157 1036 7275 1052
rect 7157 1013 7199 1036
rect 7157 979 7163 1013
rect 7197 1002 7199 1013
rect 7233 1013 7275 1036
rect 7233 1002 7235 1013
rect 7197 979 7235 1002
rect 7269 979 7275 1013
rect 7157 968 7275 979
rect 7157 940 7199 968
rect 7157 906 7163 940
rect 7197 934 7199 940
rect 7233 940 7275 968
rect 7233 934 7235 940
rect 7197 906 7235 934
rect 7269 906 7275 940
rect 7157 900 7275 906
rect 7157 867 7199 900
rect 7157 833 7163 867
rect 7197 866 7199 867
rect 7233 867 7275 900
rect 7233 866 7235 867
rect 7197 833 7235 866
rect 7269 833 7275 867
rect 7157 832 7275 833
rect 7157 798 7199 832
rect 7233 798 7275 832
rect 7157 794 7275 798
rect 7157 760 7163 794
rect 7197 764 7235 794
rect 7197 760 7199 764
rect 7157 730 7199 760
rect 7233 760 7235 764
rect 7269 760 7275 794
rect 7233 730 7275 760
rect 7157 721 7275 730
rect 7157 687 7163 721
rect 7197 696 7235 721
rect 7197 687 7199 696
rect 7157 662 7199 687
rect 7233 687 7235 696
rect 7269 687 7275 721
rect 7233 662 7275 687
rect 7157 648 7275 662
rect 7157 614 7163 648
rect 7197 628 7235 648
rect 7197 614 7199 628
rect 7157 594 7199 614
rect 7233 614 7235 628
rect 7269 614 7275 648
rect 7233 594 7275 614
rect 7157 575 7275 594
rect 7157 541 7163 575
rect 7197 560 7235 575
rect 7197 541 7199 560
rect 7157 526 7199 541
rect 7233 541 7235 560
rect 7269 541 7275 575
rect 7233 526 7275 541
rect 7157 502 7275 526
rect 7157 324 7163 502
rect 7269 364 7275 502
rect 7330 1201 7364 1213
rect 7330 1127 7364 1163
rect 11565 1201 11599 1213
rect 11565 1197 11566 1201
rect 11599 1163 11600 1167
rect 11565 1127 11600 1163
rect 11565 1123 11566 1127
rect 7330 1053 7364 1089
rect 7454 1068 7462 1102
rect 7528 1068 7530 1102
rect 7564 1068 7568 1102
rect 7632 1068 7642 1102
rect 7700 1068 7716 1102
rect 7768 1068 7790 1102
rect 7836 1068 7864 1102
rect 7904 1068 7938 1102
rect 7972 1068 8006 1102
rect 8046 1068 8074 1102
rect 8120 1068 8142 1102
rect 8194 1068 8210 1102
rect 8268 1068 8278 1102
rect 8342 1068 8346 1102
rect 8380 1068 8382 1102
rect 8448 1068 8456 1102
rect 8516 1068 8529 1102
rect 8584 1068 8602 1102
rect 8652 1068 8675 1102
rect 8720 1068 8748 1102
rect 8788 1068 8821 1102
rect 8856 1068 8890 1102
rect 8928 1068 8958 1102
rect 9001 1068 9026 1102
rect 9074 1068 9094 1102
rect 9147 1068 9162 1102
rect 9220 1068 9230 1102
rect 9293 1068 9298 1102
rect 9400 1068 9416 1102
rect 9552 1068 9564 1102
rect 9602 1068 9636 1102
rect 9671 1068 9704 1102
rect 9744 1068 9772 1102
rect 9817 1068 9840 1102
rect 9890 1068 9908 1102
rect 9963 1068 9976 1102
rect 10036 1068 10044 1102
rect 10109 1068 10112 1102
rect 10146 1068 10148 1102
rect 10214 1068 10221 1102
rect 10282 1068 10294 1102
rect 10350 1068 10367 1102
rect 10418 1068 10440 1102
rect 10486 1068 10514 1102
rect 10554 1068 10588 1102
rect 10622 1068 10656 1102
rect 10696 1068 10724 1102
rect 10770 1068 10792 1102
rect 10844 1068 10860 1102
rect 10918 1068 10928 1102
rect 10992 1068 10996 1102
rect 11030 1068 11032 1102
rect 11098 1068 11106 1102
rect 11166 1068 11180 1102
rect 11234 1068 11254 1102
rect 11302 1068 11328 1102
rect 11370 1068 11402 1102
rect 11438 1068 11472 1102
rect 11510 1068 11522 1102
rect 11599 1089 11600 1093
rect 7330 979 7364 1016
rect 11565 1053 11600 1089
rect 11565 1050 11566 1053
rect 11599 1016 11600 1019
rect 11565 979 11600 1016
rect 11565 977 11566 979
rect 7330 905 7364 943
rect 7454 912 7462 946
rect 7528 912 7530 946
rect 7564 912 7568 946
rect 7632 912 7642 946
rect 7700 912 7716 946
rect 7768 912 7790 946
rect 7836 912 7864 946
rect 7904 912 7938 946
rect 7972 912 8006 946
rect 8046 912 8074 946
rect 8120 912 8142 946
rect 8194 912 8210 946
rect 8268 912 8278 946
rect 8342 912 8346 946
rect 8380 912 8382 946
rect 8448 912 8456 946
rect 8516 912 8529 946
rect 8584 912 8602 946
rect 8652 912 8675 946
rect 8720 912 8748 946
rect 8788 912 8821 946
rect 8856 912 8890 946
rect 8928 912 8958 946
rect 9001 912 9026 946
rect 9074 912 9094 946
rect 9147 912 9162 946
rect 9220 912 9230 946
rect 9293 912 9298 946
rect 9400 912 9416 946
rect 9552 912 9564 946
rect 9602 912 9636 946
rect 9671 912 9704 946
rect 9744 912 9772 946
rect 9817 912 9840 946
rect 9890 912 9908 946
rect 9963 912 9976 946
rect 10036 912 10044 946
rect 10109 912 10112 946
rect 10146 912 10148 946
rect 10214 912 10221 946
rect 10282 912 10294 946
rect 10350 912 10367 946
rect 10418 912 10440 946
rect 10486 912 10514 946
rect 10554 912 10588 946
rect 10622 912 10656 946
rect 10696 912 10724 946
rect 10770 912 10792 946
rect 10844 912 10860 946
rect 10918 912 10928 946
rect 10992 912 10996 946
rect 11030 912 11032 946
rect 11098 912 11106 946
rect 11166 912 11180 946
rect 11234 912 11254 946
rect 11302 912 11328 946
rect 11370 912 11402 946
rect 11438 912 11472 946
rect 11510 912 11522 946
rect 11599 943 11600 945
rect 7330 831 7364 870
rect 7330 758 7364 797
rect 11565 905 11600 943
rect 11565 904 11566 905
rect 11599 870 11600 871
rect 11565 831 11600 870
rect 7454 756 7462 790
rect 7528 756 7530 790
rect 7564 756 7568 790
rect 7632 756 7642 790
rect 7700 756 7716 790
rect 7768 756 7790 790
rect 7836 756 7864 790
rect 7904 756 7938 790
rect 7972 756 8006 790
rect 8046 756 8074 790
rect 8120 756 8142 790
rect 8194 756 8210 790
rect 8268 756 8278 790
rect 8342 756 8346 790
rect 8380 756 8382 790
rect 8448 756 8456 790
rect 8516 756 8529 790
rect 8584 756 8602 790
rect 8652 756 8675 790
rect 8720 756 8748 790
rect 8788 756 8821 790
rect 8856 756 8890 790
rect 8928 756 8958 790
rect 9001 756 9026 790
rect 9074 756 9094 790
rect 9147 756 9162 790
rect 9220 756 9230 790
rect 9293 756 9298 790
rect 9400 756 9416 790
rect 9552 756 9564 790
rect 9602 756 9636 790
rect 9671 756 9704 790
rect 9744 756 9772 790
rect 9817 756 9840 790
rect 9890 756 9908 790
rect 9963 756 9976 790
rect 10036 756 10044 790
rect 10109 756 10112 790
rect 10146 756 10148 790
rect 10214 756 10221 790
rect 10282 756 10294 790
rect 10350 756 10367 790
rect 10418 756 10440 790
rect 10486 756 10514 790
rect 10554 756 10588 790
rect 10622 756 10656 790
rect 10696 756 10724 790
rect 10770 756 10792 790
rect 10844 756 10860 790
rect 10918 756 10928 790
rect 10992 756 10996 790
rect 11030 756 11032 790
rect 11098 756 11106 790
rect 11166 756 11180 790
rect 11234 756 11254 790
rect 11302 756 11328 790
rect 11370 756 11402 790
rect 11438 756 11472 790
rect 11510 756 11522 790
rect 11565 758 11600 797
rect 11599 757 11600 758
rect 7330 685 7364 723
rect 7330 612 7364 649
rect 11565 723 11566 724
rect 11565 685 11600 723
rect 11599 683 11600 685
rect 11565 649 11566 651
rect 7454 600 7462 634
rect 7528 600 7530 634
rect 7564 600 7568 634
rect 7632 600 7642 634
rect 7700 600 7716 634
rect 7768 600 7790 634
rect 7836 600 7864 634
rect 7904 600 7938 634
rect 7972 600 8006 634
rect 8046 600 8074 634
rect 8120 600 8142 634
rect 8194 600 8210 634
rect 8268 600 8278 634
rect 8342 600 8346 634
rect 8380 600 8382 634
rect 8448 600 8456 634
rect 8516 600 8529 634
rect 8584 600 8602 634
rect 8652 600 8675 634
rect 8720 600 8748 634
rect 8788 600 8821 634
rect 8856 600 8890 634
rect 8928 600 8958 634
rect 9001 600 9026 634
rect 9074 600 9094 634
rect 9147 600 9162 634
rect 9220 600 9230 634
rect 9293 600 9298 634
rect 9400 600 9416 634
rect 9552 600 9564 634
rect 9602 600 9636 634
rect 9671 600 9704 634
rect 9744 600 9772 634
rect 9817 600 9840 634
rect 9890 600 9908 634
rect 9963 600 9976 634
rect 10036 600 10044 634
rect 10109 600 10112 634
rect 10146 600 10148 634
rect 10214 600 10221 634
rect 10282 600 10294 634
rect 10350 600 10367 634
rect 10418 600 10440 634
rect 10486 600 10514 634
rect 10554 600 10588 634
rect 10622 600 10656 634
rect 10696 600 10724 634
rect 10770 600 10792 634
rect 10844 600 10860 634
rect 10918 600 10928 634
rect 10992 600 10996 634
rect 11030 600 11032 634
rect 11098 600 11106 634
rect 11166 600 11180 634
rect 11234 600 11254 634
rect 11302 600 11328 634
rect 11370 600 11402 634
rect 11438 600 11472 634
rect 11510 600 11522 634
rect 11565 612 11600 649
rect 11599 609 11600 612
rect 7330 539 7364 575
rect 7330 489 7364 501
rect 11565 575 11566 578
rect 11565 539 11600 575
rect 11599 535 11600 539
rect 11565 501 11566 505
rect 11639 1200 11645 1338
rect 11751 1200 11757 1378
rect 11639 1176 11757 1200
rect 11639 1161 11681 1176
rect 11639 1127 11645 1161
rect 11679 1142 11681 1161
rect 11715 1161 11757 1176
rect 11715 1142 11717 1161
rect 11679 1127 11717 1142
rect 11751 1127 11757 1161
rect 11639 1108 11757 1127
rect 11639 1088 11681 1108
rect 11639 1054 11645 1088
rect 11679 1074 11681 1088
rect 11715 1088 11757 1108
rect 11715 1074 11717 1088
rect 11679 1054 11717 1074
rect 11751 1054 11757 1088
rect 11639 1040 11757 1054
rect 11639 1015 11681 1040
rect 11639 981 11645 1015
rect 11679 1006 11681 1015
rect 11715 1015 11757 1040
rect 11715 1006 11717 1015
rect 11679 981 11717 1006
rect 11751 981 11757 1015
rect 11639 972 11757 981
rect 11639 942 11681 972
rect 11639 908 11645 942
rect 11679 938 11681 942
rect 11715 942 11757 972
rect 11715 938 11717 942
rect 11679 908 11717 938
rect 11751 908 11757 942
rect 11639 904 11757 908
rect 11639 870 11681 904
rect 11715 870 11757 904
rect 11639 869 11757 870
rect 11639 835 11645 869
rect 11679 836 11717 869
rect 11679 835 11681 836
rect 11639 802 11681 835
rect 11715 835 11717 836
rect 11751 835 11757 869
rect 11715 802 11757 835
rect 11639 796 11757 802
rect 11639 762 11645 796
rect 11679 768 11717 796
rect 11679 762 11681 768
rect 11639 734 11681 762
rect 11715 762 11717 768
rect 11751 762 11757 796
rect 11715 734 11757 762
rect 11639 723 11757 734
rect 11639 689 11645 723
rect 11679 700 11717 723
rect 11679 689 11681 700
rect 11639 666 11681 689
rect 11715 689 11717 700
rect 11751 689 11757 723
rect 11715 666 11757 689
rect 11639 650 11757 666
rect 11639 616 11645 650
rect 11679 632 11717 650
rect 11679 616 11681 632
rect 11639 598 11681 616
rect 11715 616 11717 632
rect 11751 616 11757 650
rect 11715 598 11757 616
rect 11639 577 11757 598
rect 11639 543 11645 577
rect 11679 564 11717 577
rect 11679 543 11681 564
rect 11639 530 11681 543
rect 11715 543 11717 564
rect 11751 543 11757 577
rect 11715 530 11757 543
rect 11639 504 11757 530
rect 11565 489 11599 501
rect 7454 444 7462 478
rect 7528 444 7530 478
rect 7564 444 7568 478
rect 7632 444 7642 478
rect 7700 444 7716 478
rect 7768 444 7790 478
rect 7836 444 7864 478
rect 7904 444 7938 478
rect 7972 444 8006 478
rect 8046 444 8074 478
rect 8120 444 8142 478
rect 8194 444 8210 478
rect 8268 444 8278 478
rect 8342 444 8346 478
rect 8380 444 8382 478
rect 8448 444 8456 478
rect 8516 444 8529 478
rect 8584 444 8602 478
rect 8652 444 8675 478
rect 8720 444 8748 478
rect 8788 444 8821 478
rect 8856 444 8890 478
rect 8928 444 8958 478
rect 9001 444 9026 478
rect 9074 444 9094 478
rect 9147 444 9162 478
rect 9220 444 9230 478
rect 9293 444 9298 478
rect 9400 444 9416 478
rect 9552 444 9564 478
rect 9602 444 9636 478
rect 9671 444 9704 478
rect 9744 444 9772 478
rect 9817 444 9840 478
rect 9890 444 9908 478
rect 9963 444 9976 478
rect 10036 444 10044 478
rect 10109 444 10112 478
rect 10146 444 10148 478
rect 10214 444 10221 478
rect 10282 444 10294 478
rect 10350 444 10367 478
rect 10418 444 10440 478
rect 10486 444 10514 478
rect 10554 444 10588 478
rect 10622 444 10656 478
rect 10696 444 10724 478
rect 10770 444 10792 478
rect 10844 444 10860 478
rect 10918 444 10928 478
rect 10992 444 10996 478
rect 11030 444 11032 478
rect 11098 444 11106 478
rect 11166 444 11180 478
rect 11234 444 11254 478
rect 11302 444 11328 478
rect 11370 444 11402 478
rect 11438 444 11472 478
rect 11510 444 11522 478
rect 11639 470 11645 504
rect 11679 496 11717 504
rect 11679 470 11681 496
rect 11639 462 11681 470
rect 11715 470 11717 496
rect 11751 470 11757 504
rect 11715 462 11757 470
rect 11639 431 11757 462
rect 11639 397 11645 431
rect 11679 428 11717 431
rect 11679 397 11681 428
rect 11639 394 11681 397
rect 11715 397 11717 428
rect 11751 397 11757 431
rect 11715 394 11757 397
rect 11639 364 11757 394
rect 7269 359 11757 364
rect 7298 358 7332 359
rect 7366 358 7400 359
rect 7434 358 7468 359
rect 7502 358 7536 359
rect 7570 358 7604 359
rect 7298 325 7308 358
rect 7366 325 7381 358
rect 7434 325 7454 358
rect 7502 325 7527 358
rect 7570 325 7600 358
rect 7638 325 7672 359
rect 7706 358 7740 359
rect 7774 358 7808 359
rect 7842 358 7876 359
rect 7910 358 7944 359
rect 7978 358 8012 359
rect 8046 358 8080 359
rect 8114 358 8148 359
rect 7707 325 7740 358
rect 7780 325 7808 358
rect 7853 325 7876 358
rect 7926 325 7944 358
rect 7999 325 8012 358
rect 8072 325 8080 358
rect 8145 325 8148 358
rect 8182 358 8216 359
rect 8250 358 8284 359
rect 8318 358 8352 359
rect 8386 358 8420 359
rect 8454 358 8488 359
rect 8522 358 8556 359
rect 8590 358 8624 359
rect 8658 358 8692 359
rect 8726 358 8760 359
rect 8794 358 8828 359
rect 8862 358 8896 359
rect 8930 358 8964 359
rect 8998 358 9032 359
rect 9066 358 9100 359
rect 9134 358 9168 359
rect 9202 358 9236 359
rect 9270 358 9304 359
rect 9338 358 9372 359
rect 9406 358 9440 359
rect 9474 358 9508 359
rect 9542 358 9576 359
rect 9610 358 9644 359
rect 9678 358 9712 359
rect 9746 358 9780 359
rect 9814 358 9848 359
rect 9882 358 9916 359
rect 9950 358 9984 359
rect 10018 358 10052 359
rect 10086 358 10120 359
rect 10154 358 10188 359
rect 10222 358 10256 359
rect 10290 358 10324 359
rect 10358 358 10392 359
rect 10426 358 10460 359
rect 10494 358 10528 359
rect 10562 358 10596 359
rect 10630 358 10664 359
rect 10698 358 10732 359
rect 10766 358 10800 359
rect 10834 358 10868 359
rect 10902 358 10936 359
rect 10970 358 11004 359
rect 11038 358 11072 359
rect 11106 358 11140 359
rect 11174 358 11208 359
rect 11242 358 11276 359
rect 11310 358 11344 359
rect 11378 358 11412 359
rect 11446 358 11480 359
rect 11514 358 11548 359
rect 11582 358 11616 359
rect 11650 358 11757 359
rect 8182 325 8184 358
rect 8250 325 8257 358
rect 8318 325 8330 358
rect 8386 325 8403 358
rect 8454 325 8476 358
rect 8522 325 8549 358
rect 7269 324 7308 325
rect 7342 324 7381 325
rect 7415 324 7454 325
rect 7488 324 7527 325
rect 7561 324 7600 325
rect 7634 324 7673 325
rect 7707 324 7746 325
rect 7780 324 7819 325
rect 7853 324 7892 325
rect 7926 324 7965 325
rect 7999 324 8038 325
rect 8072 324 8111 325
rect 8145 324 8184 325
rect 8218 324 8257 325
rect 8291 324 8330 325
rect 8364 324 8403 325
rect 8437 324 8476 325
rect 8510 324 8549 325
rect 7157 286 8549 324
rect 7157 252 7235 286
rect 7269 252 7308 286
rect 7342 252 7381 286
rect 7415 252 7454 286
rect 7488 252 7527 286
rect 7561 252 7600 286
rect 7634 252 7673 286
rect 7707 252 7746 286
rect 7780 252 7819 286
rect 7853 252 7892 286
rect 7926 252 7965 286
rect 7999 252 8038 286
rect 8072 252 8111 286
rect 8145 252 8184 286
rect 8218 252 8257 286
rect 8291 252 8330 286
rect 8364 252 8403 286
rect 8437 252 8476 286
rect 8510 252 8549 286
rect 11679 324 11717 358
rect 11751 324 11757 358
rect 11679 252 11757 324
rect 7157 246 11757 252
rect 11894 1425 12012 1463
rect 11894 1391 11900 1425
rect 11934 1391 11972 1425
rect 12006 1391 12012 1425
rect 11894 1352 12012 1391
rect 11894 1318 11900 1352
rect 11934 1318 11972 1352
rect 12006 1318 12012 1352
rect 11894 1279 12012 1318
rect 11894 1245 11900 1279
rect 11934 1245 11972 1279
rect 12006 1245 12012 1279
rect 11894 1206 12012 1245
rect 11894 1172 11900 1206
rect 11934 1172 11972 1206
rect 12006 1172 12012 1206
rect 11894 1133 12012 1172
rect 11894 1099 11900 1133
rect 11934 1099 11972 1133
rect 12006 1099 12012 1133
rect 11894 1059 12012 1099
rect 11894 1025 11900 1059
rect 11934 1025 11972 1059
rect 12006 1025 12012 1059
rect 11894 985 12012 1025
rect 11894 951 11900 985
rect 11934 951 11972 985
rect 12006 951 12012 985
rect 11894 911 12012 951
rect 11894 877 11900 911
rect 11934 877 11972 911
rect 12006 877 12012 911
rect 11894 837 12012 877
rect 11894 803 11900 837
rect 11934 803 11972 837
rect 12006 803 12012 837
rect 11894 763 12012 803
rect 11894 729 11900 763
rect 11934 729 11972 763
rect 12006 729 12012 763
rect 11894 689 12012 729
rect 11894 655 11900 689
rect 11934 655 11972 689
rect 12006 655 12012 689
rect 11894 615 12012 655
rect 11894 581 11900 615
rect 11934 581 11972 615
rect 12006 581 12012 615
rect 11894 541 12012 581
rect 11894 507 11900 541
rect 11934 507 11972 541
rect 12006 507 12012 541
rect 11894 467 12012 507
rect 11894 433 11900 467
rect 11934 433 11972 467
rect 12006 433 12012 467
rect 11894 393 12012 433
rect 11894 359 11900 393
rect 11934 359 11972 393
rect 12006 359 12012 393
rect 11894 319 12012 359
rect 11894 285 11900 319
rect 11934 285 11972 319
rect 12006 285 12012 319
rect 6876 177 6882 243
rect 2008 171 6882 177
rect 6988 177 6994 243
rect 11894 245 12012 285
rect 11894 211 11900 245
rect 11934 211 11972 245
rect 12006 211 12012 245
rect 11894 177 12012 211
rect 6988 171 12012 177
rect 167 137 206 171
rect 240 169 279 171
rect 313 169 352 171
rect 386 169 425 171
rect 459 169 498 171
rect 532 169 571 171
rect 605 169 644 171
rect 678 169 717 171
rect 751 169 790 171
rect 824 169 863 171
rect 897 169 936 171
rect 970 169 1009 171
rect 1043 169 1082 171
rect 1116 169 1155 171
rect 1189 169 1228 171
rect 1262 169 1301 171
rect 1335 169 1374 171
rect 1408 169 1447 171
rect 1481 169 1520 171
rect 1554 169 1593 171
rect 1627 169 1666 171
rect 1700 169 1739 171
rect 1773 169 1812 171
rect 1846 169 1885 171
rect 1872 137 1885 169
rect 2008 137 2031 171
rect 2065 169 2104 171
rect 2138 169 2177 171
rect 2211 169 2250 171
rect 2284 169 2323 171
rect 2357 169 2396 171
rect 2065 137 2103 169
rect 55 135 63 137
rect 165 135 206 137
rect 55 101 206 135
rect 55 99 138 101
rect 55 65 133 99
rect 172 67 206 101
rect 1872 135 1906 137
rect 2008 135 2103 137
rect 1872 101 2103 135
rect 1872 99 2035 101
rect 1872 67 1885 99
rect 167 65 206 67
rect 240 65 279 67
rect 313 65 352 67
rect 386 65 425 67
rect 459 65 498 67
rect 532 65 571 67
rect 605 65 644 67
rect 678 65 717 67
rect 751 65 790 67
rect 824 65 863 67
rect 897 65 936 67
rect 970 65 1009 67
rect 1043 65 1082 67
rect 1116 65 1155 67
rect 1189 65 1228 67
rect 1262 65 1301 67
rect 1335 65 1374 67
rect 1408 65 1447 67
rect 1481 65 1520 67
rect 1554 65 1593 67
rect 1627 65 1666 67
rect 1700 65 1739 67
rect 1773 65 1812 67
rect 1846 65 1885 67
rect 1919 65 1958 99
rect 1992 65 2031 99
rect 2069 67 2103 101
rect 11934 137 11972 171
rect 12006 137 12012 171
rect 2065 65 2104 67
rect 2138 65 2177 67
rect 2211 65 2250 67
rect 2284 65 2323 67
rect 2357 65 2396 67
rect 11934 65 12012 137
rect 55 59 12012 65
rect -462 -88 -409 -54
rect -375 -88 -322 -54
rect -288 -88 -236 -54
rect -202 -88 -150 -54
rect -496 -164 -116 -88
rect -462 -198 -409 -164
rect -375 -198 -322 -164
rect -288 -198 -236 -164
rect -202 -198 -150 -164
rect 5611 -1153 7982 -1147
rect 5611 -1187 5691 -1153
rect 5725 -1154 5765 -1153
rect 5799 -1154 5839 -1153
rect 5873 -1154 5913 -1153
rect 5947 -1154 5987 -1153
rect 6021 -1154 6062 -1153
rect 6096 -1154 6137 -1153
rect 6171 -1154 6212 -1153
rect 6246 -1154 6287 -1153
rect 6321 -1154 6397 -1153
rect 6431 -1154 6470 -1153
rect 6504 -1154 6543 -1153
rect 6577 -1154 6616 -1153
rect 5732 -1187 5765 -1154
rect 5611 -1188 5698 -1187
rect 5732 -1188 5766 -1187
rect 5800 -1188 5834 -1154
rect 5873 -1187 5902 -1154
rect 5947 -1187 5970 -1154
rect 6021 -1187 6038 -1154
rect 6096 -1187 6106 -1154
rect 6171 -1187 6174 -1154
rect 5868 -1188 5902 -1187
rect 5936 -1188 5970 -1187
rect 6004 -1188 6038 -1187
rect 6072 -1188 6106 -1187
rect 6140 -1188 6174 -1187
rect 6208 -1187 6212 -1154
rect 6276 -1187 6287 -1154
rect 6208 -1188 6242 -1187
rect 6276 -1188 6310 -1187
rect 6344 -1188 6378 -1154
rect 6431 -1187 6446 -1154
rect 6504 -1187 6514 -1154
rect 6577 -1187 6582 -1154
rect 6412 -1188 6446 -1187
rect 6480 -1188 6514 -1187
rect 6548 -1188 6582 -1187
rect 6650 -1154 6689 -1153
rect 6723 -1154 6762 -1153
rect 6796 -1154 6835 -1153
rect 6869 -1154 6908 -1153
rect 6942 -1154 6982 -1153
rect 7016 -1154 7056 -1153
rect 7090 -1154 7130 -1153
rect 7164 -1154 7204 -1153
rect 7238 -1154 7278 -1153
rect 7312 -1154 7352 -1153
rect 7386 -1154 7426 -1153
rect 7460 -1154 7500 -1153
rect 6616 -1188 6650 -1187
rect 6684 -1187 6689 -1154
rect 6752 -1187 6762 -1154
rect 6820 -1187 6835 -1154
rect 6888 -1187 6908 -1154
rect 6956 -1187 6982 -1154
rect 7024 -1187 7056 -1154
rect 6684 -1188 6718 -1187
rect 6752 -1188 6786 -1187
rect 6820 -1188 6854 -1187
rect 6888 -1188 6922 -1187
rect 6956 -1188 6990 -1187
rect 7024 -1188 7058 -1187
rect 7092 -1188 7126 -1154
rect 7164 -1187 7194 -1154
rect 7238 -1187 7262 -1154
rect 7312 -1187 7330 -1154
rect 7386 -1187 7398 -1154
rect 7460 -1187 7466 -1154
rect 7160 -1188 7194 -1187
rect 7228 -1188 7262 -1187
rect 7296 -1188 7330 -1187
rect 7364 -1188 7398 -1187
rect 7432 -1188 7466 -1187
rect 7534 -1154 7574 -1153
rect 7608 -1154 7648 -1153
rect 7682 -1154 7722 -1153
rect 7756 -1154 7796 -1153
rect 7830 -1154 7870 -1153
rect 7904 -1154 7982 -1153
rect 7500 -1188 7534 -1187
rect 7568 -1187 7574 -1154
rect 7636 -1187 7648 -1154
rect 7704 -1187 7722 -1154
rect 7772 -1187 7796 -1154
rect 7840 -1187 7870 -1154
rect 7568 -1188 7602 -1187
rect 7636 -1188 7670 -1187
rect 7704 -1188 7738 -1187
rect 7772 -1188 7806 -1187
rect 7840 -1188 7874 -1187
rect 7908 -1188 7982 -1154
rect 5611 -1193 7982 -1188
rect 5611 -1222 5657 -1193
rect 5611 -1259 5617 -1222
rect 5651 -1259 5657 -1222
rect 5611 -1290 5657 -1259
rect 7936 -1231 7982 -1193
rect 5611 -1338 5617 -1290
rect 5651 -1338 5657 -1290
rect 5850 -1304 5852 -1270
rect 5900 -1304 5927 -1270
rect 5968 -1304 6002 -1270
rect 6036 -1304 6070 -1270
rect 6111 -1304 6138 -1270
rect 6186 -1304 6206 -1270
rect 6261 -1304 6274 -1270
rect 6336 -1304 6342 -1270
rect 6376 -1304 6377 -1270
rect 6444 -1304 6452 -1270
rect 6512 -1304 6527 -1270
rect 6580 -1304 6602 -1270
rect 6648 -1304 6676 -1270
rect 6716 -1304 6750 -1270
rect 6784 -1304 6818 -1270
rect 6858 -1304 6886 -1270
rect 6932 -1304 6954 -1270
rect 7006 -1304 7022 -1270
rect 7080 -1304 7090 -1270
rect 7154 -1304 7158 -1270
rect 7192 -1304 7194 -1270
rect 7260 -1304 7268 -1270
rect 7328 -1304 7342 -1270
rect 7396 -1304 7416 -1270
rect 7464 -1304 7490 -1270
rect 7532 -1304 7564 -1270
rect 7600 -1304 7634 -1270
rect 7672 -1304 7702 -1270
rect 7746 -1304 7770 -1270
rect 7936 -1296 7942 -1231
rect 7976 -1296 7982 -1231
rect 7936 -1309 7982 -1296
rect 5611 -1358 5657 -1338
rect 5611 -1417 5617 -1358
rect 5651 -1417 5657 -1358
rect 5611 -1426 5657 -1417
rect 5611 -1460 5617 -1426
rect 5651 -1460 5657 -1426
rect 5611 -1462 5657 -1460
rect 5611 -1528 5617 -1462
rect 5651 -1528 5657 -1462
rect 5611 -1541 5657 -1528
rect 5611 -1596 5617 -1541
rect 5651 -1596 5657 -1541
rect 5611 -1620 5657 -1596
rect 5611 -1654 5617 -1620
rect 5651 -1654 5657 -1620
rect 5611 -1698 5657 -1654
rect 5611 -1758 5617 -1698
rect 5651 -1758 5657 -1698
rect 5611 -1776 5657 -1758
rect 5611 -1826 5617 -1776
rect 5651 -1826 5657 -1776
rect 5611 -1854 5657 -1826
rect 5611 -1894 5617 -1854
rect 5651 -1894 5657 -1854
rect 5734 -1327 5768 -1315
rect 5734 -1399 5768 -1365
rect 7936 -1364 7942 -1309
rect 7976 -1364 7982 -1309
rect 7936 -1387 7982 -1364
rect 5734 -1472 5768 -1436
rect 5850 -1460 5852 -1426
rect 5900 -1460 5927 -1426
rect 5968 -1460 6002 -1426
rect 6036 -1460 6070 -1426
rect 6111 -1460 6138 -1426
rect 6186 -1460 6206 -1426
rect 6261 -1460 6274 -1426
rect 6336 -1460 6342 -1426
rect 6376 -1460 6377 -1426
rect 6444 -1460 6452 -1426
rect 6512 -1460 6527 -1426
rect 6580 -1460 6602 -1426
rect 6648 -1460 6676 -1426
rect 6716 -1460 6750 -1426
rect 6784 -1460 6818 -1426
rect 6858 -1460 6886 -1426
rect 6932 -1460 6954 -1426
rect 7006 -1460 7022 -1426
rect 7080 -1460 7090 -1426
rect 7154 -1460 7158 -1426
rect 7192 -1460 7194 -1426
rect 7260 -1460 7268 -1426
rect 7328 -1460 7342 -1426
rect 7396 -1460 7416 -1426
rect 7464 -1460 7490 -1426
rect 7532 -1460 7564 -1426
rect 7600 -1460 7634 -1426
rect 7672 -1460 7702 -1426
rect 7746 -1460 7770 -1426
rect 7936 -1432 7942 -1387
rect 7976 -1432 7982 -1387
rect 5734 -1545 5768 -1507
rect 5734 -1617 5768 -1579
rect 7936 -1465 7982 -1432
rect 7936 -1500 7942 -1465
rect 7976 -1500 7982 -1465
rect 7936 -1534 7982 -1500
rect 7936 -1577 7942 -1534
rect 7976 -1577 7982 -1534
rect 5850 -1616 5852 -1582
rect 5900 -1616 5927 -1582
rect 5968 -1616 6002 -1582
rect 6036 -1616 6070 -1582
rect 6111 -1616 6138 -1582
rect 6186 -1616 6206 -1582
rect 6261 -1616 6274 -1582
rect 6336 -1616 6342 -1582
rect 6376 -1616 6377 -1582
rect 6444 -1616 6452 -1582
rect 6512 -1616 6527 -1582
rect 6580 -1616 6602 -1582
rect 6648 -1616 6676 -1582
rect 6716 -1616 6750 -1582
rect 6784 -1616 6818 -1582
rect 6858 -1616 6886 -1582
rect 6932 -1616 6954 -1582
rect 7006 -1616 7022 -1582
rect 7080 -1616 7090 -1582
rect 7154 -1616 7158 -1582
rect 7192 -1616 7194 -1582
rect 7260 -1616 7268 -1582
rect 7328 -1616 7342 -1582
rect 7396 -1616 7416 -1582
rect 7464 -1616 7490 -1582
rect 7532 -1616 7564 -1582
rect 7600 -1616 7634 -1582
rect 7672 -1616 7702 -1582
rect 7746 -1616 7770 -1582
rect 7936 -1602 7982 -1577
rect 5734 -1689 5768 -1652
rect 5734 -1761 5768 -1725
rect 7936 -1656 7942 -1602
rect 7976 -1656 7982 -1602
rect 7936 -1670 7982 -1656
rect 7936 -1735 7942 -1670
rect 7976 -1735 7982 -1670
rect 7936 -1738 7982 -1735
rect 5850 -1772 5852 -1738
rect 5900 -1772 5927 -1738
rect 5968 -1772 6002 -1738
rect 6036 -1772 6070 -1738
rect 6111 -1772 6138 -1738
rect 6186 -1772 6206 -1738
rect 6261 -1772 6274 -1738
rect 6336 -1772 6342 -1738
rect 6376 -1772 6377 -1738
rect 6444 -1772 6452 -1738
rect 6512 -1772 6527 -1738
rect 6580 -1772 6602 -1738
rect 6648 -1772 6676 -1738
rect 6716 -1772 6750 -1738
rect 6784 -1772 6818 -1738
rect 6858 -1772 6886 -1738
rect 6932 -1772 6954 -1738
rect 7006 -1772 7022 -1738
rect 7080 -1772 7090 -1738
rect 7154 -1772 7158 -1738
rect 7192 -1772 7194 -1738
rect 7260 -1772 7268 -1738
rect 7328 -1772 7342 -1738
rect 7396 -1772 7416 -1738
rect 7464 -1772 7490 -1738
rect 7532 -1772 7564 -1738
rect 7600 -1772 7634 -1738
rect 7672 -1772 7702 -1738
rect 7746 -1772 7770 -1738
rect 7936 -1772 7942 -1738
rect 7976 -1772 7982 -1738
rect 5734 -1833 5768 -1798
rect 5734 -1883 5768 -1871
rect 7936 -1780 7982 -1772
rect 7936 -1840 7942 -1780
rect 7976 -1840 7982 -1780
rect 7936 -1859 7982 -1840
rect 5611 -1928 5657 -1894
rect 5850 -1928 5852 -1894
rect 5900 -1928 5927 -1894
rect 5968 -1928 6002 -1894
rect 6036 -1928 6070 -1894
rect 6111 -1928 6138 -1894
rect 6186 -1928 6206 -1894
rect 6261 -1928 6274 -1894
rect 6336 -1928 6342 -1894
rect 6376 -1928 6377 -1894
rect 6444 -1928 6452 -1894
rect 6512 -1928 6527 -1894
rect 6580 -1928 6602 -1894
rect 6648 -1928 6676 -1894
rect 6716 -1928 6750 -1894
rect 6784 -1928 6818 -1894
rect 6858 -1928 6886 -1894
rect 6932 -1928 6954 -1894
rect 7006 -1928 7022 -1894
rect 7080 -1928 7090 -1894
rect 7154 -1928 7158 -1894
rect 7192 -1928 7194 -1894
rect 7260 -1928 7268 -1894
rect 7328 -1928 7342 -1894
rect 7396 -1928 7416 -1894
rect 7464 -1928 7490 -1894
rect 7532 -1928 7564 -1894
rect 7600 -1928 7634 -1894
rect 7672 -1928 7702 -1894
rect 7746 -1928 7770 -1894
rect 7936 -1908 7942 -1859
rect 7976 -1908 7982 -1859
rect 5611 -1966 5617 -1928
rect 5651 -1966 5657 -1928
rect 5611 -2004 5657 -1966
rect 7936 -1938 7982 -1908
rect 7936 -1976 7942 -1938
rect 7976 -1976 7982 -1938
rect 7936 -2004 7982 -1976
rect 5611 -2010 7982 -2004
rect 5611 -2044 5685 -2010
rect 5723 -2044 5753 -2010
rect 5796 -2044 5821 -2010
rect 5869 -2044 5889 -2010
rect 5942 -2044 5957 -2010
rect 6015 -2044 6025 -2010
rect 6088 -2044 6093 -2010
rect 6195 -2044 6200 -2010
rect 6263 -2044 6273 -2010
rect 6331 -2044 6346 -2010
rect 6399 -2044 6419 -2010
rect 6467 -2044 6492 -2010
rect 6535 -2044 6565 -2010
rect 6603 -2044 6637 -2010
rect 6672 -2044 6705 -2010
rect 6745 -2044 6773 -2010
rect 6818 -2044 6841 -2010
rect 6891 -2044 6909 -2010
rect 6964 -2044 6977 -2010
rect 7037 -2044 7045 -2010
rect 7110 -2044 7113 -2010
rect 7147 -2044 7149 -2010
rect 7215 -2044 7222 -2010
rect 7283 -2044 7294 -2010
rect 7351 -2044 7366 -2010
rect 7419 -2044 7438 -2010
rect 7487 -2044 7510 -2010
rect 7555 -2044 7582 -2010
rect 7623 -2044 7654 -2010
rect 7691 -2044 7725 -2010
rect 7760 -2044 7793 -2010
rect 7832 -2044 7861 -2010
rect 7904 -2044 7982 -2010
rect 5611 -2050 7982 -2044
<< viali >>
rect -496 1460 -462 1494
rect -409 1460 -375 1494
rect -322 1460 -288 1494
rect -236 1460 -202 1494
rect -150 1460 -116 1494
rect -496 1350 -462 1384
rect -409 1350 -375 1384
rect -322 1350 -288 1384
rect -236 1350 -202 1384
rect -150 1350 -116 1384
rect 61 1374 63 1408
rect 63 1374 95 1408
rect 133 1374 165 1408
rect 165 1374 167 1408
rect 61 1301 63 1335
rect 63 1301 95 1335
rect 133 1301 165 1335
rect 165 1301 167 1335
rect 61 1228 63 1262
rect 63 1228 95 1262
rect 133 1228 165 1262
rect 165 1228 167 1262
rect 61 1155 63 1189
rect 63 1155 95 1189
rect 133 1155 165 1189
rect 165 1155 167 1189
rect 61 1082 63 1116
rect 63 1082 95 1116
rect 133 1082 165 1116
rect 165 1082 167 1116
rect 61 1009 63 1043
rect 63 1009 95 1043
rect 133 1009 165 1043
rect 165 1009 167 1043
rect 61 936 63 970
rect 63 936 95 970
rect 133 936 165 970
rect 165 936 167 970
rect 61 863 63 897
rect 63 863 95 897
rect 133 863 165 897
rect 165 863 167 897
rect 61 790 63 824
rect 63 790 95 824
rect 133 790 165 824
rect 165 790 167 824
rect -497 726 -463 760
rect -410 726 -376 760
rect -323 726 -289 760
rect -236 726 -202 760
rect -150 726 -116 760
rect -497 648 -463 682
rect -410 648 -376 682
rect -323 648 -289 682
rect -236 648 -202 682
rect -150 648 -116 682
rect -497 570 -463 604
rect -410 570 -376 604
rect -323 570 -289 604
rect -236 570 -202 604
rect -150 570 -116 604
rect 61 717 63 751
rect 63 717 95 751
rect 133 717 165 751
rect 165 717 167 751
rect 61 644 63 678
rect 63 644 95 678
rect 133 644 165 678
rect 165 644 167 678
rect 61 571 63 605
rect 63 571 95 605
rect 133 571 165 605
rect 165 571 167 605
rect 61 498 63 532
rect 63 498 95 532
rect 133 498 165 532
rect 165 498 167 532
rect 61 137 63 459
rect 63 137 165 459
rect 165 137 167 459
rect 402 1392 436 1426
rect 480 1392 514 1426
rect 558 1392 592 1426
rect 636 1392 670 1426
rect 714 1392 748 1426
rect 792 1392 826 1426
rect 870 1392 904 1426
rect 949 1392 983 1426
rect 324 1320 358 1354
rect 396 1320 430 1354
rect 480 1351 514 1354
rect 558 1351 592 1354
rect 636 1351 670 1354
rect 714 1351 748 1354
rect 792 1351 826 1354
rect 870 1351 904 1354
rect 949 1351 983 1354
rect 1059 1351 1597 1426
rect 1636 1392 1670 1426
rect 1636 1351 1670 1354
rect 480 1320 492 1351
rect 492 1320 514 1351
rect 558 1320 560 1351
rect 560 1320 592 1351
rect 636 1320 662 1351
rect 662 1320 670 1351
rect 714 1320 730 1351
rect 730 1320 748 1351
rect 792 1320 798 1351
rect 798 1320 826 1351
rect 870 1320 900 1351
rect 900 1320 904 1351
rect 949 1320 968 1351
rect 968 1320 983 1351
rect 1059 1320 1131 1351
rect 1131 1320 1165 1351
rect 1165 1320 1199 1351
rect 1199 1320 1233 1351
rect 1233 1320 1267 1351
rect 1267 1320 1301 1351
rect 1301 1320 1335 1351
rect 1335 1320 1369 1351
rect 1369 1320 1403 1351
rect 1403 1320 1437 1351
rect 1437 1320 1471 1351
rect 1471 1320 1505 1351
rect 1505 1320 1539 1351
rect 1539 1320 1573 1351
rect 1573 1320 1597 1351
rect 1636 1320 1641 1351
rect 1641 1320 1670 1351
rect 1708 1316 1742 1350
rect 324 1243 358 1277
rect 396 1243 430 1277
rect 324 1166 358 1200
rect 396 1166 430 1200
rect 324 1089 358 1123
rect 396 1089 430 1123
rect 324 1012 358 1046
rect 396 1012 430 1046
rect 324 935 358 969
rect 396 935 430 969
rect 324 858 358 892
rect 396 858 430 892
rect 324 782 358 816
rect 396 782 430 816
rect 324 706 358 740
rect 396 706 430 740
rect 324 630 358 664
rect 396 630 430 664
rect 324 554 358 588
rect 396 554 430 588
rect 324 478 358 512
rect 396 478 430 512
rect 1636 1240 1670 1274
rect 1708 1240 1742 1274
rect 566 1232 600 1235
rect 641 1232 675 1235
rect 716 1232 750 1235
rect 791 1232 825 1235
rect 866 1232 900 1235
rect 940 1232 974 1235
rect 1014 1232 1048 1235
rect 1088 1232 1122 1235
rect 1162 1232 1196 1235
rect 1236 1232 1270 1235
rect 1310 1232 1344 1235
rect 1384 1232 1418 1235
rect 1458 1232 1492 1235
rect 566 1201 570 1232
rect 570 1201 600 1232
rect 641 1201 672 1232
rect 672 1201 675 1232
rect 716 1201 740 1232
rect 740 1201 750 1232
rect 791 1201 808 1232
rect 808 1201 825 1232
rect 866 1201 876 1232
rect 876 1201 900 1232
rect 940 1201 944 1232
rect 944 1201 974 1232
rect 1014 1201 1046 1232
rect 1046 1201 1048 1232
rect 1088 1201 1114 1232
rect 1114 1201 1122 1232
rect 1162 1201 1182 1232
rect 1182 1201 1196 1232
rect 1236 1201 1250 1232
rect 1250 1201 1270 1232
rect 1310 1201 1318 1232
rect 1318 1201 1344 1232
rect 1384 1201 1386 1232
rect 1386 1201 1418 1232
rect 1458 1201 1488 1232
rect 1488 1201 1492 1232
rect 476 1160 510 1175
rect 476 1141 510 1160
rect 476 1090 510 1102
rect 476 1068 510 1090
rect 1636 1164 1670 1198
rect 1708 1164 1742 1198
rect 1636 1088 1670 1122
rect 1124 1042 1148 1076
rect 1148 1042 1158 1076
rect 1202 1042 1216 1076
rect 1216 1042 1236 1076
rect 1280 1042 1284 1076
rect 1284 1042 1314 1076
rect 1358 1042 1386 1076
rect 1386 1042 1392 1076
rect 1435 1042 1454 1076
rect 1454 1042 1469 1076
rect 1512 1042 1546 1076
rect 1708 1088 1742 1122
rect 476 1020 510 1029
rect 476 995 510 1020
rect 476 950 510 956
rect 476 922 510 950
rect 1636 1012 1670 1046
rect 1708 1012 1742 1046
rect 1636 936 1670 970
rect 1708 936 1742 970
rect 566 920 600 921
rect 641 920 675 921
rect 716 920 750 921
rect 791 920 825 921
rect 866 920 900 921
rect 940 920 974 921
rect 1014 920 1048 921
rect 1088 920 1122 921
rect 1162 920 1196 921
rect 1236 920 1270 921
rect 1310 920 1344 921
rect 1384 920 1418 921
rect 1458 920 1492 921
rect 566 887 570 920
rect 570 887 600 920
rect 641 887 672 920
rect 672 887 675 920
rect 716 887 740 920
rect 740 887 750 920
rect 791 887 808 920
rect 808 887 825 920
rect 866 887 876 920
rect 876 887 900 920
rect 940 887 944 920
rect 944 887 974 920
rect 1014 887 1046 920
rect 1046 887 1048 920
rect 1088 887 1114 920
rect 1114 887 1122 920
rect 1162 887 1182 920
rect 1182 887 1196 920
rect 1236 887 1250 920
rect 1250 887 1270 920
rect 1310 887 1318 920
rect 1318 887 1344 920
rect 1384 887 1386 920
rect 1386 887 1418 920
rect 1458 887 1488 920
rect 1488 887 1492 920
rect 476 880 510 883
rect 476 849 510 880
rect 476 776 510 810
rect 1636 860 1670 894
rect 1708 860 1742 894
rect 566 756 570 790
rect 570 756 600 790
rect 641 756 672 790
rect 672 756 675 790
rect 716 756 740 790
rect 740 756 750 790
rect 791 756 808 790
rect 808 756 825 790
rect 866 756 876 790
rect 876 756 900 790
rect 940 756 944 790
rect 944 756 974 790
rect 1014 756 1046 790
rect 1046 756 1048 790
rect 1088 756 1114 790
rect 1114 756 1122 790
rect 1162 756 1182 790
rect 1182 756 1196 790
rect 1236 756 1250 790
rect 1250 756 1270 790
rect 1310 756 1318 790
rect 1318 756 1344 790
rect 1384 756 1386 790
rect 1386 756 1418 790
rect 1458 756 1488 790
rect 1488 756 1492 790
rect 1636 784 1670 818
rect 1708 784 1742 818
rect 476 706 510 738
rect 476 704 510 706
rect 476 635 510 666
rect 476 632 510 635
rect 1636 707 1670 741
rect 1708 707 1742 741
rect 1123 600 1148 634
rect 1148 600 1157 634
rect 1201 600 1216 634
rect 1216 600 1235 634
rect 1279 600 1284 634
rect 1284 600 1313 634
rect 1357 600 1386 634
rect 1386 600 1391 634
rect 1435 600 1454 634
rect 1454 600 1469 634
rect 1512 600 1546 634
rect 1636 630 1670 664
rect 1708 630 1742 664
rect 476 564 510 594
rect 476 560 510 564
rect 476 488 510 522
rect 1636 553 1670 587
rect 1708 553 1742 587
rect 566 444 570 478
rect 570 444 600 478
rect 641 444 672 478
rect 672 444 675 478
rect 716 444 740 478
rect 740 444 750 478
rect 791 444 808 478
rect 808 444 825 478
rect 866 444 876 478
rect 876 444 900 478
rect 940 444 944 478
rect 944 444 974 478
rect 1014 444 1046 478
rect 1046 444 1048 478
rect 1088 444 1114 478
rect 1114 444 1122 478
rect 1162 444 1182 478
rect 1182 444 1196 478
rect 1236 444 1250 478
rect 1250 444 1270 478
rect 1310 444 1318 478
rect 1318 444 1344 478
rect 1384 444 1386 478
rect 1386 444 1418 478
rect 1458 444 1488 478
rect 1488 444 1492 478
rect 1636 476 1670 510
rect 1708 476 1742 510
rect 324 402 358 436
rect 396 402 430 436
rect 1636 399 1670 433
rect 1708 399 1742 433
rect 324 326 358 360
rect 396 325 425 356
rect 425 325 430 356
rect 469 325 493 356
rect 493 325 503 356
rect 542 325 561 356
rect 561 325 576 356
rect 615 325 629 356
rect 629 325 649 356
rect 688 325 697 356
rect 697 325 722 356
rect 761 325 765 356
rect 765 325 795 356
rect 834 325 867 356
rect 867 325 868 356
rect 907 325 935 356
rect 935 325 941 356
rect 980 325 1003 356
rect 1003 325 1014 356
rect 1053 325 1071 356
rect 1071 325 1087 356
rect 1126 325 1139 356
rect 1139 325 1160 356
rect 1199 325 1207 356
rect 1207 325 1233 356
rect 1272 325 1275 356
rect 1275 325 1306 356
rect 1345 325 1377 356
rect 1377 325 1379 356
rect 1418 325 1445 356
rect 1445 325 1452 356
rect 1491 325 1513 356
rect 1513 325 1525 356
rect 1564 325 1581 356
rect 1581 325 1615 356
rect 1615 325 1670 356
rect 396 322 430 325
rect 469 322 503 325
rect 542 322 576 325
rect 615 322 649 325
rect 688 322 722 325
rect 761 322 795 325
rect 834 322 868 325
rect 907 322 941 325
rect 980 322 1014 325
rect 1053 322 1087 325
rect 1126 322 1160 325
rect 1199 322 1233 325
rect 1272 322 1306 325
rect 1345 322 1379 325
rect 1418 322 1452 325
rect 1491 322 1525 325
rect 396 250 430 284
rect 469 250 503 284
rect 542 250 576 284
rect 615 250 649 284
rect 688 250 722 284
rect 761 250 795 284
rect 834 250 868 284
rect 907 250 941 284
rect 980 250 1014 284
rect 1053 250 1087 284
rect 1126 250 1160 284
rect 1199 250 1233 284
rect 1272 250 1306 284
rect 1345 250 1379 284
rect 1418 250 1452 284
rect 1491 250 1525 284
rect 1564 250 1670 325
rect 1708 322 1742 356
rect 1904 1400 1906 1434
rect 1906 1400 1938 1434
rect 1976 1400 2008 1434
rect 2008 1400 2010 1434
rect 1904 1325 1906 1359
rect 1906 1325 1938 1359
rect 1976 1325 2008 1359
rect 2008 1325 2010 1359
rect 1904 1250 1906 1284
rect 1906 1250 1938 1284
rect 1976 1250 2008 1284
rect 2008 1250 2010 1284
rect 1904 1175 1906 1209
rect 1906 1175 1938 1209
rect 1976 1175 2008 1209
rect 2008 1175 2010 1209
rect 1904 1100 1906 1134
rect 1906 1100 1938 1134
rect 1976 1100 2008 1134
rect 2008 1100 2010 1134
rect 1904 1025 1906 1059
rect 1906 1025 1938 1059
rect 1976 1025 2008 1059
rect 2008 1025 2010 1059
rect 1904 950 1906 984
rect 1906 950 1938 984
rect 1976 950 2008 984
rect 2008 950 2010 984
rect 1904 875 1906 909
rect 1906 875 1938 909
rect 1976 875 2008 909
rect 2008 875 2010 909
rect 1904 801 1906 835
rect 1906 801 1938 835
rect 1976 801 2008 835
rect 2008 801 2010 835
rect 1904 727 1906 761
rect 1906 727 1938 761
rect 1976 727 2008 761
rect 2008 727 2010 761
rect 1904 653 1906 687
rect 1906 653 1938 687
rect 1976 653 2008 687
rect 2008 653 2010 687
rect 1904 579 1906 613
rect 1906 579 1938 613
rect 1976 579 2008 613
rect 2008 579 2010 613
rect 1904 505 1906 539
rect 1906 505 1938 539
rect 1976 505 2008 539
rect 2008 505 2010 539
rect 1904 431 1906 465
rect 1906 431 1938 465
rect 1976 431 2008 465
rect 2008 431 2010 465
rect 1904 357 1906 391
rect 1906 357 1938 391
rect 1976 357 2008 391
rect 2008 357 2010 391
rect 1904 283 1906 317
rect 1906 283 1938 317
rect 1976 283 2008 317
rect 2008 283 2010 317
rect 2237 1416 2271 1450
rect 2315 1416 2349 1450
rect 2393 1416 2427 1450
rect 2471 1416 2505 1450
rect 2549 1416 2583 1450
rect 2627 1416 2661 1450
rect 2705 1416 2739 1450
rect 2784 1416 2818 1450
rect 2894 1416 2928 1450
rect 2967 1416 3001 1450
rect 3040 1416 3074 1450
rect 3113 1416 3147 1450
rect 3186 1416 3220 1450
rect 3259 1416 3293 1450
rect 3332 1416 3366 1450
rect 3405 1416 3439 1450
rect 3478 1416 3512 1450
rect 3551 1416 3585 1450
rect 3624 1416 3658 1450
rect 3697 1416 3731 1450
rect 3770 1416 3804 1450
rect 3843 1416 3877 1450
rect 3916 1416 3950 1450
rect 3989 1416 4023 1450
rect 4062 1416 4096 1450
rect 4135 1416 4169 1450
rect 4208 1416 4242 1450
rect 4281 1416 4315 1450
rect 4354 1416 4388 1450
rect 4427 1416 4461 1450
rect 4500 1416 4534 1450
rect 4573 1416 4607 1450
rect 4646 1416 4680 1450
rect 4719 1416 4753 1450
rect 4792 1416 4826 1450
rect 4865 1416 4899 1450
rect 4938 1416 4972 1450
rect 5011 1416 5045 1450
rect 5084 1416 5118 1450
rect 5157 1416 5191 1450
rect 5230 1416 5264 1450
rect 5303 1416 5337 1450
rect 5376 1416 5410 1450
rect 5449 1416 5483 1450
rect 5522 1416 5556 1450
rect 5595 1416 5629 1450
rect 5668 1416 5702 1450
rect 5741 1416 5775 1450
rect 5814 1416 5848 1450
rect 5887 1416 5921 1450
rect 5961 1416 5995 1450
rect 6035 1416 6069 1450
rect 6109 1416 6143 1450
rect 6183 1416 6217 1450
rect 6257 1416 6291 1450
rect 6331 1416 6365 1450
rect 6405 1416 6439 1450
rect 6479 1416 6513 1450
rect 6553 1416 6587 1450
rect 6627 1416 6661 1450
rect 2159 1344 2193 1378
rect 2231 1344 2265 1378
rect 2315 1377 2349 1378
rect 2393 1377 2427 1378
rect 2471 1377 2505 1378
rect 2549 1377 2583 1378
rect 2627 1377 2661 1378
rect 2705 1377 2739 1378
rect 2784 1377 2818 1378
rect 2894 1377 2928 1378
rect 2967 1377 3001 1378
rect 3040 1377 3074 1378
rect 3113 1377 3147 1378
rect 3186 1377 3220 1378
rect 3259 1377 3293 1378
rect 3332 1377 3366 1378
rect 3405 1377 3439 1378
rect 3478 1377 3512 1378
rect 3551 1377 3585 1378
rect 3624 1377 3658 1378
rect 3697 1377 3731 1378
rect 3770 1377 3804 1378
rect 3843 1377 3877 1378
rect 3916 1377 3950 1378
rect 3989 1377 4023 1378
rect 4062 1377 4096 1378
rect 4135 1377 4169 1378
rect 4208 1377 4242 1378
rect 4281 1377 4315 1378
rect 4354 1377 4388 1378
rect 4427 1377 4461 1378
rect 2315 1344 2321 1377
rect 2321 1344 2349 1377
rect 2393 1344 2423 1377
rect 2423 1344 2427 1377
rect 2471 1344 2491 1377
rect 2491 1344 2505 1377
rect 2549 1344 2559 1377
rect 2559 1344 2583 1377
rect 2627 1344 2661 1377
rect 2705 1344 2729 1377
rect 2729 1344 2739 1377
rect 2784 1344 2797 1377
rect 2797 1344 2818 1377
rect 2894 1344 2899 1377
rect 2899 1344 2928 1377
rect 2967 1344 3001 1377
rect 3040 1344 3069 1377
rect 3069 1344 3074 1377
rect 3113 1344 3137 1377
rect 3137 1344 3147 1377
rect 3186 1344 3205 1377
rect 3205 1344 3220 1377
rect 3259 1344 3273 1377
rect 3273 1344 3293 1377
rect 3332 1344 3341 1377
rect 3341 1344 3366 1377
rect 3405 1344 3409 1377
rect 3409 1344 3439 1377
rect 3478 1344 3511 1377
rect 3511 1344 3512 1377
rect 3551 1344 3579 1377
rect 3579 1344 3585 1377
rect 3624 1344 3647 1377
rect 3647 1344 3658 1377
rect 3697 1344 3715 1377
rect 3715 1344 3731 1377
rect 3770 1344 3783 1377
rect 3783 1344 3804 1377
rect 3843 1344 3851 1377
rect 3851 1344 3877 1377
rect 3916 1344 3919 1377
rect 3919 1344 3950 1377
rect 3989 1344 4021 1377
rect 4021 1344 4023 1377
rect 4062 1344 4089 1377
rect 4089 1344 4096 1377
rect 4135 1344 4157 1377
rect 4157 1344 4169 1377
rect 4208 1344 4225 1377
rect 4225 1344 4242 1377
rect 4281 1344 4293 1377
rect 4293 1344 4315 1377
rect 4354 1344 4361 1377
rect 4361 1344 4388 1377
rect 4427 1344 4429 1377
rect 4429 1344 4461 1377
rect 4500 1344 4534 1378
rect 4573 1377 4607 1378
rect 4646 1377 4680 1378
rect 4719 1377 4753 1378
rect 4792 1377 4826 1378
rect 4865 1377 4899 1378
rect 4938 1377 4972 1378
rect 5011 1377 5045 1378
rect 5084 1377 5118 1378
rect 5157 1377 5191 1378
rect 5230 1377 5264 1378
rect 5303 1377 5337 1378
rect 5376 1377 5410 1378
rect 5449 1377 5483 1378
rect 5522 1377 5556 1378
rect 5595 1377 5629 1378
rect 5668 1377 5702 1378
rect 5741 1377 5775 1378
rect 5814 1377 5848 1378
rect 5887 1377 5921 1378
rect 5961 1377 5995 1378
rect 6035 1377 6069 1378
rect 6109 1377 6143 1378
rect 6183 1377 6217 1378
rect 6257 1377 6291 1378
rect 6331 1377 6365 1378
rect 6405 1377 6439 1378
rect 6479 1377 6513 1378
rect 6553 1377 6587 1378
rect 6627 1377 6733 1378
rect 4573 1344 4592 1377
rect 4592 1344 4607 1377
rect 4646 1344 4660 1377
rect 4660 1344 4680 1377
rect 4719 1344 4728 1377
rect 4728 1344 4753 1377
rect 4792 1344 4796 1377
rect 4796 1344 4826 1377
rect 4865 1344 4898 1377
rect 4898 1344 4899 1377
rect 4938 1344 4966 1377
rect 4966 1344 4972 1377
rect 5011 1344 5034 1377
rect 5034 1344 5045 1377
rect 5084 1344 5102 1377
rect 5102 1344 5118 1377
rect 5157 1344 5170 1377
rect 5170 1344 5191 1377
rect 5230 1344 5238 1377
rect 5238 1344 5264 1377
rect 5303 1344 5306 1377
rect 5306 1344 5337 1377
rect 5376 1344 5408 1377
rect 5408 1344 5410 1377
rect 5449 1344 5476 1377
rect 5476 1344 5483 1377
rect 5522 1344 5544 1377
rect 5544 1344 5556 1377
rect 5595 1344 5612 1377
rect 5612 1344 5629 1377
rect 5668 1344 5680 1377
rect 5680 1344 5702 1377
rect 5741 1344 5748 1377
rect 5748 1344 5775 1377
rect 5814 1344 5816 1377
rect 5816 1344 5848 1377
rect 5887 1344 5918 1377
rect 5918 1344 5921 1377
rect 5961 1344 5986 1377
rect 5986 1344 5995 1377
rect 6035 1344 6054 1377
rect 6054 1344 6069 1377
rect 6109 1344 6122 1377
rect 6122 1344 6143 1377
rect 6183 1344 6190 1377
rect 6190 1344 6217 1377
rect 6257 1344 6258 1377
rect 6258 1344 6291 1377
rect 6331 1344 6360 1377
rect 6360 1344 6365 1377
rect 6405 1344 6428 1377
rect 6428 1344 6439 1377
rect 6479 1344 6496 1377
rect 6496 1344 6513 1377
rect 6553 1344 6564 1377
rect 6564 1344 6587 1377
rect 6627 1343 6632 1377
rect 6632 1343 6733 1377
rect 2159 1271 2193 1305
rect 2231 1271 2265 1305
rect 2159 1198 2193 1232
rect 2231 1198 2265 1232
rect 2401 1224 2405 1258
rect 2405 1224 2435 1258
rect 2475 1224 2507 1258
rect 2507 1224 2509 1258
rect 2549 1224 2575 1258
rect 2575 1224 2583 1258
rect 2623 1224 2643 1258
rect 2643 1224 2657 1258
rect 2697 1224 2711 1258
rect 2711 1224 2731 1258
rect 2771 1224 2779 1258
rect 2779 1224 2805 1258
rect 2845 1224 2847 1258
rect 2847 1224 2879 1258
rect 2919 1224 2949 1258
rect 2949 1224 2953 1258
rect 2993 1224 3017 1258
rect 3017 1224 3027 1258
rect 3067 1224 3085 1258
rect 3085 1224 3101 1258
rect 3141 1224 3153 1258
rect 3153 1224 3175 1258
rect 3215 1224 3221 1258
rect 3221 1224 3249 1258
rect 3289 1224 3323 1258
rect 3363 1224 3391 1258
rect 3391 1224 3397 1258
rect 3437 1224 3459 1258
rect 3459 1224 3471 1258
rect 3510 1224 3527 1258
rect 3527 1224 3544 1258
rect 3583 1224 3595 1258
rect 3595 1224 3617 1258
rect 3656 1224 3663 1258
rect 3663 1224 3690 1258
rect 3729 1224 3731 1258
rect 3731 1224 3763 1258
rect 3802 1224 3833 1258
rect 3833 1224 3836 1258
rect 3875 1224 3901 1258
rect 3901 1224 3909 1258
rect 3948 1224 3969 1258
rect 3969 1224 3982 1258
rect 4021 1224 4037 1258
rect 4037 1224 4055 1258
rect 4094 1224 4105 1258
rect 4105 1224 4128 1258
rect 4167 1224 4173 1258
rect 4173 1224 4201 1258
rect 4240 1224 4241 1258
rect 4241 1224 4274 1258
rect 4313 1224 4343 1258
rect 4343 1224 4347 1258
rect 4545 1224 4549 1258
rect 4549 1224 4579 1258
rect 4618 1224 4651 1258
rect 4651 1224 4652 1258
rect 4691 1224 4719 1258
rect 4719 1224 4725 1258
rect 4764 1224 4787 1258
rect 4787 1224 4798 1258
rect 4837 1224 4855 1258
rect 4855 1224 4871 1258
rect 4910 1224 4923 1258
rect 4923 1224 4944 1258
rect 4983 1224 4991 1258
rect 4991 1224 5017 1258
rect 5056 1224 5059 1258
rect 5059 1224 5090 1258
rect 5129 1224 5161 1258
rect 5161 1224 5163 1258
rect 5202 1224 5229 1258
rect 5229 1224 5236 1258
rect 5275 1224 5297 1258
rect 5297 1224 5309 1258
rect 5348 1224 5365 1258
rect 5365 1224 5382 1258
rect 5421 1224 5433 1258
rect 5433 1224 5455 1258
rect 5495 1224 5501 1258
rect 5501 1224 5529 1258
rect 5569 1224 5603 1258
rect 5643 1224 5671 1258
rect 5671 1224 5677 1258
rect 5717 1224 5739 1258
rect 5739 1224 5751 1258
rect 5791 1224 5807 1258
rect 5807 1224 5825 1258
rect 5865 1224 5875 1258
rect 5875 1224 5899 1258
rect 5939 1224 5943 1258
rect 5943 1224 5973 1258
rect 6013 1224 6045 1258
rect 6045 1224 6047 1258
rect 6087 1224 6113 1258
rect 6113 1224 6121 1258
rect 6161 1224 6181 1258
rect 6181 1224 6195 1258
rect 6235 1224 6249 1258
rect 6249 1224 6269 1258
rect 6309 1224 6317 1258
rect 6317 1224 6343 1258
rect 6383 1224 6385 1258
rect 6385 1224 6417 1258
rect 6457 1224 6487 1258
rect 6487 1224 6491 1258
rect 2159 1125 2193 1159
rect 2231 1125 2265 1159
rect 2159 1052 2193 1086
rect 2231 1052 2265 1086
rect 2159 979 2193 1013
rect 2231 979 2265 1013
rect 2159 906 2193 940
rect 2231 906 2265 940
rect 2159 833 2193 867
rect 2231 833 2265 867
rect 2159 760 2193 794
rect 2231 760 2265 794
rect 2159 687 2193 721
rect 2231 687 2265 721
rect 2159 614 2193 648
rect 2231 614 2265 648
rect 2159 541 2193 575
rect 2231 541 2265 575
rect 2311 1197 2345 1201
rect 2311 1167 2345 1197
rect 2311 1123 2345 1128
rect 2311 1094 2345 1123
rect 6547 1197 6581 1201
rect 6547 1167 6581 1197
rect 6547 1123 6581 1129
rect 2401 1068 2405 1102
rect 2405 1068 2435 1102
rect 2475 1068 2507 1102
rect 2507 1068 2509 1102
rect 2549 1068 2575 1102
rect 2575 1068 2583 1102
rect 2623 1068 2643 1102
rect 2643 1068 2657 1102
rect 2697 1068 2711 1102
rect 2711 1068 2731 1102
rect 2771 1068 2779 1102
rect 2779 1068 2805 1102
rect 2845 1068 2847 1102
rect 2847 1068 2879 1102
rect 2919 1068 2949 1102
rect 2949 1068 2953 1102
rect 2993 1068 3017 1102
rect 3017 1068 3027 1102
rect 3067 1068 3085 1102
rect 3085 1068 3101 1102
rect 3141 1068 3153 1102
rect 3153 1068 3175 1102
rect 3215 1068 3221 1102
rect 3221 1068 3249 1102
rect 3289 1068 3323 1102
rect 3363 1068 3391 1102
rect 3391 1068 3397 1102
rect 3437 1068 3459 1102
rect 3459 1068 3471 1102
rect 3510 1068 3527 1102
rect 3527 1068 3544 1102
rect 3583 1068 3595 1102
rect 3595 1068 3617 1102
rect 3656 1068 3663 1102
rect 3663 1068 3690 1102
rect 3729 1068 3731 1102
rect 3731 1068 3763 1102
rect 3802 1068 3833 1102
rect 3833 1068 3836 1102
rect 3875 1068 3901 1102
rect 3901 1068 3909 1102
rect 3948 1068 3969 1102
rect 3969 1068 3982 1102
rect 4021 1068 4037 1102
rect 4037 1068 4055 1102
rect 4094 1068 4105 1102
rect 4105 1068 4128 1102
rect 4167 1068 4173 1102
rect 4173 1068 4201 1102
rect 4240 1068 4241 1102
rect 4241 1068 4274 1102
rect 4313 1068 4343 1102
rect 4343 1068 4347 1102
rect 4545 1068 4549 1102
rect 4549 1068 4579 1102
rect 4618 1068 4651 1102
rect 4651 1068 4652 1102
rect 4691 1068 4719 1102
rect 4719 1068 4725 1102
rect 4764 1068 4787 1102
rect 4787 1068 4798 1102
rect 4837 1068 4855 1102
rect 4855 1068 4871 1102
rect 4910 1068 4923 1102
rect 4923 1068 4944 1102
rect 4983 1068 4991 1102
rect 4991 1068 5017 1102
rect 5056 1068 5059 1102
rect 5059 1068 5090 1102
rect 5129 1068 5161 1102
rect 5161 1068 5163 1102
rect 5202 1068 5229 1102
rect 5229 1068 5236 1102
rect 5275 1068 5297 1102
rect 5297 1068 5309 1102
rect 5348 1068 5365 1102
rect 5365 1068 5382 1102
rect 5421 1068 5433 1102
rect 5433 1068 5455 1102
rect 5495 1068 5501 1102
rect 5501 1068 5529 1102
rect 5569 1068 5603 1102
rect 5643 1068 5671 1102
rect 5671 1068 5677 1102
rect 5717 1068 5739 1102
rect 5739 1068 5751 1102
rect 5791 1068 5807 1102
rect 5807 1068 5825 1102
rect 5865 1068 5875 1102
rect 5875 1068 5899 1102
rect 5939 1068 5943 1102
rect 5943 1068 5973 1102
rect 6013 1068 6045 1102
rect 6045 1068 6047 1102
rect 6087 1068 6113 1102
rect 6113 1068 6121 1102
rect 6161 1068 6181 1102
rect 6181 1068 6195 1102
rect 6235 1068 6249 1102
rect 6249 1068 6269 1102
rect 6309 1068 6317 1102
rect 6317 1068 6343 1102
rect 6383 1068 6385 1102
rect 6385 1068 6417 1102
rect 6457 1068 6487 1102
rect 6487 1068 6491 1102
rect 6547 1095 6581 1123
rect 2311 1049 2345 1055
rect 2311 1021 2345 1049
rect 2311 974 2345 981
rect 2311 947 2345 974
rect 6547 1049 6581 1056
rect 6547 1022 6581 1049
rect 6547 974 6581 983
rect 6547 949 6581 974
rect 2401 912 2405 946
rect 2405 912 2435 946
rect 2475 912 2507 946
rect 2507 912 2509 946
rect 2549 912 2575 946
rect 2575 912 2583 946
rect 2623 912 2643 946
rect 2643 912 2657 946
rect 2697 912 2711 946
rect 2711 912 2731 946
rect 2771 912 2779 946
rect 2779 912 2805 946
rect 2845 912 2847 946
rect 2847 912 2879 946
rect 2919 912 2949 946
rect 2949 912 2953 946
rect 2993 912 3017 946
rect 3017 912 3027 946
rect 3067 912 3085 946
rect 3085 912 3101 946
rect 3141 912 3153 946
rect 3153 912 3175 946
rect 3215 912 3221 946
rect 3221 912 3249 946
rect 3289 912 3323 946
rect 3363 912 3391 946
rect 3391 912 3397 946
rect 3437 912 3459 946
rect 3459 912 3471 946
rect 3510 912 3527 946
rect 3527 912 3544 946
rect 3583 912 3595 946
rect 3595 912 3617 946
rect 3656 912 3663 946
rect 3663 912 3690 946
rect 3729 912 3731 946
rect 3731 912 3763 946
rect 3802 912 3833 946
rect 3833 912 3836 946
rect 3875 912 3901 946
rect 3901 912 3909 946
rect 3948 912 3969 946
rect 3969 912 3982 946
rect 4021 912 4037 946
rect 4037 912 4055 946
rect 4094 912 4105 946
rect 4105 912 4128 946
rect 4167 912 4173 946
rect 4173 912 4201 946
rect 4240 912 4241 946
rect 4241 912 4274 946
rect 4313 912 4343 946
rect 4343 912 4347 946
rect 4545 912 4549 946
rect 4549 912 4579 946
rect 4618 912 4651 946
rect 4651 912 4652 946
rect 4691 912 4719 946
rect 4719 912 4725 946
rect 4764 912 4787 946
rect 4787 912 4798 946
rect 4837 912 4855 946
rect 4855 912 4871 946
rect 4910 912 4923 946
rect 4923 912 4944 946
rect 4983 912 4991 946
rect 4991 912 5017 946
rect 5056 912 5059 946
rect 5059 912 5090 946
rect 5129 912 5161 946
rect 5161 912 5163 946
rect 5202 912 5229 946
rect 5229 912 5236 946
rect 5275 912 5297 946
rect 5297 912 5309 946
rect 5348 912 5365 946
rect 5365 912 5382 946
rect 5421 912 5433 946
rect 5433 912 5455 946
rect 5495 912 5501 946
rect 5501 912 5529 946
rect 5569 912 5603 946
rect 5643 912 5671 946
rect 5671 912 5677 946
rect 5717 912 5739 946
rect 5739 912 5751 946
rect 5791 912 5807 946
rect 5807 912 5825 946
rect 5865 912 5875 946
rect 5875 912 5899 946
rect 5939 912 5943 946
rect 5943 912 5973 946
rect 6013 912 6045 946
rect 6045 912 6047 946
rect 6087 912 6113 946
rect 6113 912 6121 946
rect 6161 912 6181 946
rect 6181 912 6195 946
rect 6235 912 6249 946
rect 6249 912 6269 946
rect 6309 912 6317 946
rect 6317 912 6343 946
rect 6383 912 6385 946
rect 6385 912 6417 946
rect 6457 912 6487 946
rect 6487 912 6491 946
rect 2311 899 2345 907
rect 2311 873 2345 899
rect 2311 824 2345 833
rect 2311 799 2345 824
rect 6547 899 6581 910
rect 6547 876 6581 899
rect 6547 824 6581 837
rect 6547 803 6581 824
rect 2311 749 2345 759
rect 2401 756 2405 790
rect 2405 756 2435 790
rect 2475 756 2507 790
rect 2507 756 2509 790
rect 2549 756 2575 790
rect 2575 756 2583 790
rect 2623 756 2643 790
rect 2643 756 2657 790
rect 2697 756 2711 790
rect 2711 756 2731 790
rect 2771 756 2779 790
rect 2779 756 2805 790
rect 2845 756 2847 790
rect 2847 756 2879 790
rect 2919 756 2949 790
rect 2949 756 2953 790
rect 2993 756 3017 790
rect 3017 756 3027 790
rect 3067 756 3085 790
rect 3085 756 3101 790
rect 3141 756 3153 790
rect 3153 756 3175 790
rect 3215 756 3221 790
rect 3221 756 3249 790
rect 3289 756 3323 790
rect 3363 756 3391 790
rect 3391 756 3397 790
rect 3437 756 3459 790
rect 3459 756 3471 790
rect 3510 756 3527 790
rect 3527 756 3544 790
rect 3583 756 3595 790
rect 3595 756 3617 790
rect 3656 756 3663 790
rect 3663 756 3690 790
rect 3729 756 3731 790
rect 3731 756 3763 790
rect 3802 756 3833 790
rect 3833 756 3836 790
rect 3875 756 3901 790
rect 3901 756 3909 790
rect 3948 756 3969 790
rect 3969 756 3982 790
rect 4021 756 4037 790
rect 4037 756 4055 790
rect 4094 756 4105 790
rect 4105 756 4128 790
rect 4167 756 4173 790
rect 4173 756 4201 790
rect 4240 756 4241 790
rect 4241 756 4274 790
rect 4313 756 4343 790
rect 4343 756 4347 790
rect 4545 756 4549 790
rect 4549 756 4579 790
rect 4618 756 4651 790
rect 4651 756 4652 790
rect 4691 756 4719 790
rect 4719 756 4725 790
rect 4764 756 4787 790
rect 4787 756 4798 790
rect 4837 756 4855 790
rect 4855 756 4871 790
rect 4910 756 4923 790
rect 4923 756 4944 790
rect 4983 756 4991 790
rect 4991 756 5017 790
rect 5056 756 5059 790
rect 5059 756 5090 790
rect 5129 756 5161 790
rect 5161 756 5163 790
rect 5202 756 5229 790
rect 5229 756 5236 790
rect 5275 756 5297 790
rect 5297 756 5309 790
rect 5348 756 5365 790
rect 5365 756 5382 790
rect 5421 756 5433 790
rect 5433 756 5455 790
rect 5495 756 5501 790
rect 5501 756 5529 790
rect 5569 756 5603 790
rect 5643 756 5671 790
rect 5671 756 5677 790
rect 5717 756 5739 790
rect 5739 756 5751 790
rect 5791 756 5807 790
rect 5807 756 5825 790
rect 5865 756 5875 790
rect 5875 756 5899 790
rect 5939 756 5943 790
rect 5943 756 5973 790
rect 6013 756 6045 790
rect 6045 756 6047 790
rect 6087 756 6113 790
rect 6113 756 6121 790
rect 6161 756 6181 790
rect 6181 756 6195 790
rect 6235 756 6249 790
rect 6249 756 6269 790
rect 6309 756 6317 790
rect 6317 756 6343 790
rect 6383 756 6385 790
rect 6385 756 6417 790
rect 6457 756 6487 790
rect 6487 756 6491 790
rect 2311 725 2345 749
rect 2311 674 2345 685
rect 2311 651 2345 674
rect 6547 749 6581 764
rect 6547 730 6581 749
rect 6547 674 6581 691
rect 6547 657 6581 674
rect 2401 600 2405 634
rect 2405 600 2435 634
rect 2475 600 2507 634
rect 2507 600 2509 634
rect 2549 600 2575 634
rect 2575 600 2583 634
rect 2623 600 2643 634
rect 2643 600 2657 634
rect 2697 600 2711 634
rect 2711 600 2731 634
rect 2771 600 2779 634
rect 2779 600 2805 634
rect 2845 600 2847 634
rect 2847 600 2879 634
rect 2919 600 2949 634
rect 2949 600 2953 634
rect 2993 600 3017 634
rect 3017 600 3027 634
rect 3067 600 3085 634
rect 3085 600 3101 634
rect 3141 600 3153 634
rect 3153 600 3175 634
rect 3215 600 3221 634
rect 3221 600 3249 634
rect 3289 600 3323 634
rect 3363 600 3391 634
rect 3391 600 3397 634
rect 3437 600 3459 634
rect 3459 600 3471 634
rect 3510 600 3527 634
rect 3527 600 3544 634
rect 3583 600 3595 634
rect 3595 600 3617 634
rect 3656 600 3663 634
rect 3663 600 3690 634
rect 3729 600 3731 634
rect 3731 600 3763 634
rect 3802 600 3833 634
rect 3833 600 3836 634
rect 3875 600 3901 634
rect 3901 600 3909 634
rect 3948 600 3969 634
rect 3969 600 3982 634
rect 4021 600 4037 634
rect 4037 600 4055 634
rect 4094 600 4105 634
rect 4105 600 4128 634
rect 4167 600 4173 634
rect 4173 600 4201 634
rect 4240 600 4241 634
rect 4241 600 4274 634
rect 4313 600 4343 634
rect 4343 600 4347 634
rect 4545 600 4549 634
rect 4549 600 4579 634
rect 4618 600 4651 634
rect 4651 600 4652 634
rect 4691 600 4719 634
rect 4719 600 4725 634
rect 4764 600 4787 634
rect 4787 600 4798 634
rect 4837 600 4855 634
rect 4855 600 4871 634
rect 4910 600 4923 634
rect 4923 600 4944 634
rect 4983 600 4991 634
rect 4991 600 5017 634
rect 5056 600 5059 634
rect 5059 600 5090 634
rect 5129 600 5161 634
rect 5161 600 5163 634
rect 5202 600 5229 634
rect 5229 600 5236 634
rect 5275 600 5297 634
rect 5297 600 5309 634
rect 5348 600 5365 634
rect 5365 600 5382 634
rect 5421 600 5433 634
rect 5433 600 5455 634
rect 5495 600 5501 634
rect 5501 600 5529 634
rect 5569 600 5603 634
rect 5643 600 5671 634
rect 5671 600 5677 634
rect 5717 600 5739 634
rect 5739 600 5751 634
rect 5791 600 5807 634
rect 5807 600 5825 634
rect 5865 600 5875 634
rect 5875 600 5899 634
rect 5939 600 5943 634
rect 5943 600 5973 634
rect 6013 600 6045 634
rect 6045 600 6047 634
rect 6087 600 6113 634
rect 6113 600 6121 634
rect 6161 600 6181 634
rect 6181 600 6195 634
rect 6235 600 6249 634
rect 6249 600 6269 634
rect 6309 600 6317 634
rect 6317 600 6343 634
rect 6383 600 6385 634
rect 6385 600 6417 634
rect 6457 600 6487 634
rect 6487 600 6491 634
rect 6627 1308 6733 1343
rect 6627 1274 6663 1308
rect 6663 1274 6697 1308
rect 6697 1274 6733 1308
rect 6627 1240 6733 1274
rect 6627 1206 6663 1240
rect 6663 1206 6697 1240
rect 6697 1206 6733 1240
rect 6627 1200 6733 1206
rect 6627 1127 6661 1161
rect 6699 1127 6733 1161
rect 6627 1054 6661 1088
rect 6699 1054 6733 1088
rect 6627 981 6661 1015
rect 6699 981 6733 1015
rect 6627 908 6661 942
rect 6699 908 6733 942
rect 6627 835 6661 869
rect 6699 835 6733 869
rect 6627 762 6661 796
rect 6699 762 6733 796
rect 6627 689 6661 723
rect 6699 689 6733 723
rect 6627 616 6661 650
rect 6699 616 6733 650
rect 2159 496 2265 502
rect 2159 462 2195 496
rect 2195 462 2229 496
rect 2229 462 2265 496
rect 2159 428 2265 462
rect 2159 394 2195 428
rect 2195 394 2229 428
rect 2229 394 2265 428
rect 2159 359 2265 394
rect 6627 543 6661 577
rect 6699 543 6733 577
rect 2401 444 2405 478
rect 2405 444 2435 478
rect 2475 444 2507 478
rect 2507 444 2509 478
rect 2549 444 2575 478
rect 2575 444 2583 478
rect 2623 444 2643 478
rect 2643 444 2657 478
rect 2697 444 2711 478
rect 2711 444 2731 478
rect 2771 444 2779 478
rect 2779 444 2805 478
rect 2845 444 2847 478
rect 2847 444 2879 478
rect 2919 444 2949 478
rect 2949 444 2953 478
rect 2993 444 3017 478
rect 3017 444 3027 478
rect 3067 444 3085 478
rect 3085 444 3101 478
rect 3141 444 3153 478
rect 3153 444 3175 478
rect 3215 444 3221 478
rect 3221 444 3249 478
rect 3289 444 3323 478
rect 3363 444 3391 478
rect 3391 444 3397 478
rect 3437 444 3459 478
rect 3459 444 3471 478
rect 3510 444 3527 478
rect 3527 444 3544 478
rect 3583 444 3595 478
rect 3595 444 3617 478
rect 3656 444 3663 478
rect 3663 444 3690 478
rect 3729 444 3731 478
rect 3731 444 3763 478
rect 3802 444 3833 478
rect 3833 444 3836 478
rect 3875 444 3901 478
rect 3901 444 3909 478
rect 3948 444 3969 478
rect 3969 444 3982 478
rect 4021 444 4037 478
rect 4037 444 4055 478
rect 4094 444 4105 478
rect 4105 444 4128 478
rect 4167 444 4173 478
rect 4173 444 4201 478
rect 4240 444 4241 478
rect 4241 444 4274 478
rect 4313 444 4343 478
rect 4343 444 4347 478
rect 4545 444 4549 478
rect 4549 444 4579 478
rect 4618 444 4651 478
rect 4651 444 4652 478
rect 4691 444 4719 478
rect 4719 444 4725 478
rect 4764 444 4787 478
rect 4787 444 4798 478
rect 4837 444 4855 478
rect 4855 444 4871 478
rect 4910 444 4923 478
rect 4923 444 4944 478
rect 4983 444 4991 478
rect 4991 444 5017 478
rect 5056 444 5059 478
rect 5059 444 5090 478
rect 5129 444 5161 478
rect 5161 444 5163 478
rect 5202 444 5229 478
rect 5229 444 5236 478
rect 5275 444 5297 478
rect 5297 444 5309 478
rect 5348 444 5365 478
rect 5365 444 5382 478
rect 5421 444 5433 478
rect 5433 444 5455 478
rect 5495 444 5501 478
rect 5501 444 5529 478
rect 5569 444 5603 478
rect 5643 444 5671 478
rect 5671 444 5677 478
rect 5717 444 5739 478
rect 5739 444 5751 478
rect 5791 444 5807 478
rect 5807 444 5825 478
rect 5865 444 5875 478
rect 5875 444 5899 478
rect 5939 444 5943 478
rect 5943 444 5973 478
rect 6013 444 6045 478
rect 6045 444 6047 478
rect 6087 444 6113 478
rect 6113 444 6121 478
rect 6161 444 6181 478
rect 6181 444 6195 478
rect 6235 444 6249 478
rect 6249 444 6269 478
rect 6309 444 6317 478
rect 6317 444 6343 478
rect 6383 444 6385 478
rect 6385 444 6417 478
rect 6457 444 6487 478
rect 6487 444 6491 478
rect 6627 470 6661 504
rect 6699 470 6733 504
rect 6627 397 6661 431
rect 6699 397 6733 431
rect 2159 325 2260 359
rect 2260 325 2265 359
rect 2304 325 2328 358
rect 2328 325 2338 358
rect 2377 325 2396 358
rect 2396 325 2411 358
rect 2450 325 2464 358
rect 2464 325 2484 358
rect 2523 325 2532 358
rect 2532 325 2566 358
rect 2566 325 2600 358
rect 2600 325 2634 358
rect 2634 325 2668 358
rect 2668 325 2702 358
rect 2702 325 2736 358
rect 2736 325 2770 358
rect 2770 325 2804 358
rect 2804 325 2838 358
rect 2838 325 2872 358
rect 2872 325 2906 358
rect 2906 325 2940 358
rect 2940 325 2974 358
rect 2974 325 3008 358
rect 3008 325 3042 358
rect 3042 325 3076 358
rect 3076 325 3110 358
rect 3110 325 3144 358
rect 3144 325 3178 358
rect 3178 325 3212 358
rect 3212 325 3246 358
rect 3246 325 3280 358
rect 3280 325 3314 358
rect 3314 325 3348 358
rect 3348 325 3382 358
rect 3382 325 3416 358
rect 3416 325 3450 358
rect 3450 325 3484 358
rect 3484 325 3518 358
rect 3518 325 3552 358
rect 3552 325 3586 358
rect 3586 325 3620 358
rect 3620 325 3654 358
rect 3654 325 3688 358
rect 3688 325 3722 358
rect 3722 325 3756 358
rect 3756 325 3790 358
rect 3790 325 3824 358
rect 3824 325 3858 358
rect 3858 325 3892 358
rect 3892 325 3926 358
rect 3926 325 3960 358
rect 3960 325 3994 358
rect 3994 325 4028 358
rect 4028 325 4062 358
rect 4062 325 4096 358
rect 4096 325 4130 358
rect 4130 325 4164 358
rect 4164 325 4198 358
rect 4198 325 4232 358
rect 4232 325 4266 358
rect 4266 325 4300 358
rect 4300 325 4334 358
rect 4334 325 4368 358
rect 4368 325 4402 358
rect 4402 325 4436 358
rect 4436 325 4470 358
rect 4470 325 4504 358
rect 4504 325 4538 358
rect 4538 325 4572 358
rect 4572 325 4606 358
rect 4606 325 4640 358
rect 4640 325 4674 358
rect 4674 325 4708 358
rect 4708 325 4742 358
rect 4742 325 4776 358
rect 4776 325 4810 358
rect 4810 325 4844 358
rect 4844 325 4878 358
rect 4878 325 4912 358
rect 4912 325 4946 358
rect 4946 325 4980 358
rect 4980 325 5014 358
rect 5014 325 5048 358
rect 5048 325 5082 358
rect 5082 325 5116 358
rect 5116 325 5150 358
rect 5150 325 5184 358
rect 5184 325 5218 358
rect 5218 325 5252 358
rect 5252 325 5286 358
rect 5286 325 5320 358
rect 5320 325 5354 358
rect 5354 325 5388 358
rect 5388 325 5422 358
rect 5422 325 5456 358
rect 5456 325 5490 358
rect 5490 325 5524 358
rect 5524 325 5558 358
rect 5558 325 5592 358
rect 5592 325 5626 358
rect 5626 325 5660 358
rect 5660 325 5694 358
rect 5694 325 5728 358
rect 5728 325 5762 358
rect 5762 325 5796 358
rect 5796 325 5830 358
rect 5830 325 5864 358
rect 5864 325 5898 358
rect 5898 325 5932 358
rect 5932 325 5966 358
rect 5966 325 6000 358
rect 6000 325 6034 358
rect 6034 325 6068 358
rect 6068 325 6102 358
rect 6102 325 6136 358
rect 6136 325 6170 358
rect 6170 325 6204 358
rect 6204 325 6238 358
rect 6238 325 6272 358
rect 6272 325 6306 358
rect 6306 325 6340 358
rect 6340 325 6374 358
rect 6374 325 6408 358
rect 6408 325 6442 358
rect 6442 325 6476 358
rect 6476 325 6510 358
rect 6510 325 6544 358
rect 6544 325 6578 358
rect 6578 325 6661 358
rect 2159 324 2265 325
rect 2304 324 2338 325
rect 2377 324 2411 325
rect 2450 324 2484 325
rect 2231 252 2265 286
rect 2304 252 2338 286
rect 2377 252 2411 286
rect 2450 252 2484 286
rect 2523 252 6661 325
rect 6699 324 6733 358
rect 6882 1382 6884 1416
rect 6884 1382 6916 1416
rect 6954 1382 6986 1416
rect 6986 1382 6988 1416
rect 6882 1309 6884 1343
rect 6884 1309 6916 1343
rect 6954 1309 6986 1343
rect 6986 1309 6988 1343
rect 6882 1236 6884 1270
rect 6884 1236 6916 1270
rect 6954 1236 6986 1270
rect 6986 1236 6988 1270
rect 6882 1163 6884 1197
rect 6884 1163 6916 1197
rect 6954 1163 6986 1197
rect 6986 1163 6988 1197
rect 6882 1090 6884 1124
rect 6884 1090 6916 1124
rect 6954 1090 6986 1124
rect 6986 1090 6988 1124
rect 6882 1017 6884 1051
rect 6884 1017 6916 1051
rect 6954 1017 6986 1051
rect 6986 1017 6988 1051
rect 6882 944 6884 978
rect 6884 944 6916 978
rect 6954 944 6986 978
rect 6986 944 6988 978
rect 6882 871 6884 905
rect 6884 871 6916 905
rect 6954 871 6986 905
rect 6986 871 6988 905
rect 6882 798 6884 832
rect 6884 798 6916 832
rect 6954 798 6986 832
rect 6986 798 6988 832
rect 6882 725 6884 759
rect 6884 725 6916 759
rect 6954 725 6986 759
rect 6986 725 6988 759
rect 6882 652 6884 686
rect 6884 652 6916 686
rect 6954 652 6986 686
rect 6986 652 6988 686
rect 6882 579 6884 613
rect 6884 579 6916 613
rect 6954 579 6986 613
rect 6986 579 6988 613
rect 6882 505 6884 539
rect 6884 505 6916 539
rect 6954 505 6986 539
rect 6986 505 6988 539
rect 6882 431 6884 465
rect 6884 431 6916 465
rect 6954 431 6986 465
rect 6986 431 6988 465
rect 6882 357 6884 391
rect 6884 357 6916 391
rect 6954 357 6986 391
rect 6986 357 6988 391
rect 6882 283 6884 317
rect 6884 283 6916 317
rect 6954 283 6986 317
rect 6986 283 6988 317
rect 1904 209 1906 243
rect 1906 209 1938 243
rect 1976 209 2008 243
rect 2008 209 2010 243
rect 7241 1416 7275 1450
rect 7319 1416 7353 1450
rect 7397 1416 7431 1450
rect 7475 1416 7509 1450
rect 7553 1416 7587 1450
rect 7631 1416 7665 1450
rect 7709 1416 7743 1450
rect 7788 1416 7822 1450
rect 7163 1344 7197 1378
rect 7235 1377 7269 1378
rect 7319 1377 7353 1378
rect 7397 1377 7431 1378
rect 7475 1377 7509 1378
rect 7553 1377 7587 1378
rect 7631 1377 7665 1378
rect 7709 1377 7743 1378
rect 7788 1377 7822 1378
rect 7898 1377 11460 1450
rect 11499 1416 11533 1450
rect 11572 1416 11606 1450
rect 11645 1416 11679 1450
rect 11499 1377 11533 1378
rect 11572 1377 11606 1378
rect 7235 1344 7264 1377
rect 7264 1344 7269 1377
rect 7319 1344 7332 1377
rect 7332 1344 7353 1377
rect 7397 1344 7400 1377
rect 7400 1344 7431 1377
rect 7475 1344 7502 1377
rect 7502 1344 7509 1377
rect 7553 1344 7570 1377
rect 7570 1344 7587 1377
rect 7631 1344 7638 1377
rect 7638 1344 7665 1377
rect 7709 1344 7740 1377
rect 7740 1344 7743 1377
rect 7788 1344 7808 1377
rect 7808 1344 7822 1377
rect 7898 1344 7910 1377
rect 7910 1344 7944 1377
rect 7944 1344 7978 1377
rect 7978 1344 8012 1377
rect 8012 1344 8046 1377
rect 8046 1344 8080 1377
rect 8080 1344 8114 1377
rect 8114 1344 8148 1377
rect 8148 1344 8182 1377
rect 8182 1344 8216 1377
rect 8216 1344 8250 1377
rect 8250 1344 8284 1377
rect 8284 1344 8318 1377
rect 8318 1344 8352 1377
rect 8352 1344 8386 1377
rect 8386 1344 8420 1377
rect 8420 1344 8454 1377
rect 8454 1344 8488 1377
rect 8488 1344 8522 1377
rect 8522 1344 8556 1377
rect 8556 1344 8590 1377
rect 8590 1344 8624 1377
rect 8624 1344 8658 1377
rect 8658 1344 8692 1377
rect 8692 1344 8726 1377
rect 8726 1344 8760 1377
rect 8760 1344 8794 1377
rect 8794 1344 8828 1377
rect 8828 1344 8862 1377
rect 8862 1344 8896 1377
rect 8896 1344 8930 1377
rect 8930 1344 8964 1377
rect 8964 1344 8998 1377
rect 8998 1344 9032 1377
rect 9032 1344 9066 1377
rect 9066 1344 9100 1377
rect 9100 1344 9134 1377
rect 9134 1344 9168 1377
rect 9168 1344 9202 1377
rect 9202 1344 9236 1377
rect 9236 1344 9270 1377
rect 9270 1344 9304 1377
rect 9304 1344 9338 1377
rect 9338 1344 9372 1377
rect 9372 1344 9406 1377
rect 9406 1344 9500 1377
rect 9500 1344 9534 1377
rect 9534 1344 9568 1377
rect 9568 1344 9602 1377
rect 9602 1344 9636 1377
rect 9636 1344 9670 1377
rect 9670 1344 9704 1377
rect 9704 1344 9738 1377
rect 9738 1344 9772 1377
rect 9772 1344 9806 1377
rect 9806 1344 9840 1377
rect 9840 1344 9874 1377
rect 9874 1344 9908 1377
rect 9908 1344 9942 1377
rect 9942 1344 9976 1377
rect 9976 1344 10010 1377
rect 10010 1344 10044 1377
rect 10044 1344 10078 1377
rect 10078 1344 10112 1377
rect 10112 1344 10146 1377
rect 10146 1344 10180 1377
rect 10180 1344 10214 1377
rect 10214 1344 10248 1377
rect 10248 1344 10282 1377
rect 10282 1344 10316 1377
rect 10316 1344 10350 1377
rect 10350 1344 10384 1377
rect 10384 1344 10418 1377
rect 10418 1344 10452 1377
rect 10452 1344 10486 1377
rect 10486 1344 10520 1377
rect 10520 1344 10554 1377
rect 10554 1344 10588 1377
rect 10588 1344 10622 1377
rect 10622 1344 10656 1377
rect 10656 1344 10690 1377
rect 10690 1344 10724 1377
rect 10724 1344 10758 1377
rect 10758 1344 10792 1377
rect 10792 1344 10826 1377
rect 10826 1344 10860 1377
rect 10860 1344 10894 1377
rect 10894 1344 10928 1377
rect 10928 1344 10962 1377
rect 10962 1344 10996 1377
rect 10996 1344 11030 1377
rect 11030 1344 11064 1377
rect 11064 1344 11098 1377
rect 11098 1344 11132 1377
rect 11132 1344 11166 1377
rect 11166 1344 11200 1377
rect 11200 1344 11234 1377
rect 11234 1344 11268 1377
rect 11268 1344 11302 1377
rect 11302 1344 11336 1377
rect 11336 1344 11370 1377
rect 11370 1344 11404 1377
rect 11404 1344 11438 1377
rect 11438 1344 11460 1377
rect 11499 1344 11506 1377
rect 11506 1344 11533 1377
rect 11572 1344 11574 1377
rect 11574 1344 11606 1377
rect 7163 1271 7197 1305
rect 7235 1271 7269 1305
rect 7163 1198 7197 1232
rect 7235 1198 7269 1232
rect 7420 1224 7454 1258
rect 7494 1224 7496 1258
rect 7496 1224 7528 1258
rect 7568 1224 7598 1258
rect 7598 1224 7602 1258
rect 7642 1224 7666 1258
rect 7666 1224 7676 1258
rect 7716 1224 7734 1258
rect 7734 1224 7750 1258
rect 7790 1224 7802 1258
rect 7802 1224 7824 1258
rect 7864 1224 7870 1258
rect 7870 1224 7898 1258
rect 7938 1224 7972 1258
rect 8012 1224 8040 1258
rect 8040 1224 8046 1258
rect 8086 1224 8108 1258
rect 8108 1224 8120 1258
rect 8160 1224 8176 1258
rect 8176 1224 8194 1258
rect 8234 1224 8244 1258
rect 8244 1224 8268 1258
rect 8308 1224 8312 1258
rect 8312 1224 8342 1258
rect 8382 1224 8414 1258
rect 8414 1224 8416 1258
rect 8456 1224 8482 1258
rect 8482 1224 8490 1258
rect 8529 1224 8550 1258
rect 8550 1224 8563 1258
rect 8602 1224 8618 1258
rect 8618 1224 8636 1258
rect 8675 1224 8686 1258
rect 8686 1224 8709 1258
rect 8748 1224 8754 1258
rect 8754 1224 8782 1258
rect 8821 1224 8822 1258
rect 8822 1224 8855 1258
rect 8894 1224 8924 1258
rect 8924 1224 8928 1258
rect 8967 1224 8992 1258
rect 8992 1224 9001 1258
rect 9040 1224 9060 1258
rect 9060 1224 9074 1258
rect 9113 1224 9128 1258
rect 9128 1224 9147 1258
rect 9186 1224 9196 1258
rect 9196 1224 9220 1258
rect 9259 1224 9264 1258
rect 9264 1224 9293 1258
rect 9332 1224 9366 1258
rect 9564 1224 9568 1258
rect 9568 1224 9598 1258
rect 9637 1224 9670 1258
rect 9670 1224 9671 1258
rect 9710 1224 9738 1258
rect 9738 1224 9744 1258
rect 9783 1224 9806 1258
rect 9806 1224 9817 1258
rect 9856 1224 9874 1258
rect 9874 1224 9890 1258
rect 9929 1224 9942 1258
rect 9942 1224 9963 1258
rect 10002 1224 10010 1258
rect 10010 1224 10036 1258
rect 10075 1224 10078 1258
rect 10078 1224 10109 1258
rect 10148 1224 10180 1258
rect 10180 1224 10182 1258
rect 10221 1224 10248 1258
rect 10248 1224 10255 1258
rect 10294 1224 10316 1258
rect 10316 1224 10328 1258
rect 10367 1224 10384 1258
rect 10384 1224 10401 1258
rect 10440 1224 10452 1258
rect 10452 1224 10474 1258
rect 10514 1224 10520 1258
rect 10520 1224 10548 1258
rect 10588 1224 10622 1258
rect 10662 1224 10690 1258
rect 10690 1224 10696 1258
rect 10736 1224 10758 1258
rect 10758 1224 10770 1258
rect 10810 1224 10826 1258
rect 10826 1224 10844 1258
rect 10884 1224 10894 1258
rect 10894 1224 10918 1258
rect 10958 1224 10962 1258
rect 10962 1224 10992 1258
rect 11032 1224 11064 1258
rect 11064 1224 11066 1258
rect 11106 1224 11132 1258
rect 11132 1224 11140 1258
rect 11180 1224 11200 1258
rect 11200 1224 11214 1258
rect 11254 1224 11268 1258
rect 11268 1224 11288 1258
rect 11328 1224 11336 1258
rect 11336 1224 11362 1258
rect 11402 1224 11404 1258
rect 11404 1224 11436 1258
rect 11476 1224 11506 1258
rect 11506 1224 11510 1258
rect 7163 1125 7197 1159
rect 7235 1125 7269 1159
rect 7163 1052 7197 1086
rect 7235 1052 7269 1086
rect 7163 979 7197 1013
rect 7235 979 7269 1013
rect 7163 906 7197 940
rect 7235 906 7269 940
rect 7163 833 7197 867
rect 7235 833 7269 867
rect 7163 760 7197 794
rect 7235 760 7269 794
rect 7163 687 7197 721
rect 7235 687 7269 721
rect 7163 614 7197 648
rect 7235 614 7269 648
rect 7163 541 7197 575
rect 7235 541 7269 575
rect 7163 492 7269 502
rect 7163 458 7199 492
rect 7199 458 7233 492
rect 7233 458 7269 492
rect 7163 424 7269 458
rect 7163 390 7199 424
rect 7199 390 7233 424
rect 7233 390 7269 424
rect 7163 359 7269 390
rect 7330 1197 7364 1201
rect 7330 1167 7364 1197
rect 7330 1123 7364 1127
rect 7330 1093 7364 1123
rect 11566 1197 11600 1201
rect 11566 1167 11599 1197
rect 11599 1167 11600 1197
rect 11566 1123 11600 1127
rect 7420 1068 7454 1102
rect 7494 1068 7496 1102
rect 7496 1068 7528 1102
rect 7568 1068 7598 1102
rect 7598 1068 7602 1102
rect 7642 1068 7666 1102
rect 7666 1068 7676 1102
rect 7716 1068 7734 1102
rect 7734 1068 7750 1102
rect 7790 1068 7802 1102
rect 7802 1068 7824 1102
rect 7864 1068 7870 1102
rect 7870 1068 7898 1102
rect 7938 1068 7972 1102
rect 8012 1068 8040 1102
rect 8040 1068 8046 1102
rect 8086 1068 8108 1102
rect 8108 1068 8120 1102
rect 8160 1068 8176 1102
rect 8176 1068 8194 1102
rect 8234 1068 8244 1102
rect 8244 1068 8268 1102
rect 8308 1068 8312 1102
rect 8312 1068 8342 1102
rect 8382 1068 8414 1102
rect 8414 1068 8416 1102
rect 8456 1068 8482 1102
rect 8482 1068 8490 1102
rect 8529 1068 8550 1102
rect 8550 1068 8563 1102
rect 8602 1068 8618 1102
rect 8618 1068 8636 1102
rect 8675 1068 8686 1102
rect 8686 1068 8709 1102
rect 8748 1068 8754 1102
rect 8754 1068 8782 1102
rect 8821 1068 8822 1102
rect 8822 1068 8855 1102
rect 8894 1068 8924 1102
rect 8924 1068 8928 1102
rect 8967 1068 8992 1102
rect 8992 1068 9001 1102
rect 9040 1068 9060 1102
rect 9060 1068 9074 1102
rect 9113 1068 9128 1102
rect 9128 1068 9147 1102
rect 9186 1068 9196 1102
rect 9196 1068 9220 1102
rect 9259 1068 9264 1102
rect 9264 1068 9293 1102
rect 9332 1068 9366 1102
rect 9564 1068 9568 1102
rect 9568 1068 9598 1102
rect 9637 1068 9670 1102
rect 9670 1068 9671 1102
rect 9710 1068 9738 1102
rect 9738 1068 9744 1102
rect 9783 1068 9806 1102
rect 9806 1068 9817 1102
rect 9856 1068 9874 1102
rect 9874 1068 9890 1102
rect 9929 1068 9942 1102
rect 9942 1068 9963 1102
rect 10002 1068 10010 1102
rect 10010 1068 10036 1102
rect 10075 1068 10078 1102
rect 10078 1068 10109 1102
rect 10148 1068 10180 1102
rect 10180 1068 10182 1102
rect 10221 1068 10248 1102
rect 10248 1068 10255 1102
rect 10294 1068 10316 1102
rect 10316 1068 10328 1102
rect 10367 1068 10384 1102
rect 10384 1068 10401 1102
rect 10440 1068 10452 1102
rect 10452 1068 10474 1102
rect 10514 1068 10520 1102
rect 10520 1068 10548 1102
rect 10588 1068 10622 1102
rect 10662 1068 10690 1102
rect 10690 1068 10696 1102
rect 10736 1068 10758 1102
rect 10758 1068 10770 1102
rect 10810 1068 10826 1102
rect 10826 1068 10844 1102
rect 10884 1068 10894 1102
rect 10894 1068 10918 1102
rect 10958 1068 10962 1102
rect 10962 1068 10992 1102
rect 11032 1068 11064 1102
rect 11064 1068 11066 1102
rect 11106 1068 11132 1102
rect 11132 1068 11140 1102
rect 11180 1068 11200 1102
rect 11200 1068 11214 1102
rect 11254 1068 11268 1102
rect 11268 1068 11288 1102
rect 11328 1068 11336 1102
rect 11336 1068 11362 1102
rect 11402 1068 11404 1102
rect 11404 1068 11436 1102
rect 11476 1068 11506 1102
rect 11506 1068 11510 1102
rect 11566 1093 11599 1123
rect 11599 1093 11600 1123
rect 7330 1050 7364 1053
rect 7330 1019 7364 1050
rect 7330 977 7364 979
rect 7330 945 7364 977
rect 11566 1050 11600 1053
rect 11566 1019 11599 1050
rect 11599 1019 11600 1050
rect 11566 977 11600 979
rect 7420 912 7454 946
rect 7494 912 7496 946
rect 7496 912 7528 946
rect 7568 912 7598 946
rect 7598 912 7602 946
rect 7642 912 7666 946
rect 7666 912 7676 946
rect 7716 912 7734 946
rect 7734 912 7750 946
rect 7790 912 7802 946
rect 7802 912 7824 946
rect 7864 912 7870 946
rect 7870 912 7898 946
rect 7938 912 7972 946
rect 8012 912 8040 946
rect 8040 912 8046 946
rect 8086 912 8108 946
rect 8108 912 8120 946
rect 8160 912 8176 946
rect 8176 912 8194 946
rect 8234 912 8244 946
rect 8244 912 8268 946
rect 8308 912 8312 946
rect 8312 912 8342 946
rect 8382 912 8414 946
rect 8414 912 8416 946
rect 8456 912 8482 946
rect 8482 912 8490 946
rect 8529 912 8550 946
rect 8550 912 8563 946
rect 8602 912 8618 946
rect 8618 912 8636 946
rect 8675 912 8686 946
rect 8686 912 8709 946
rect 8748 912 8754 946
rect 8754 912 8782 946
rect 8821 912 8822 946
rect 8822 912 8855 946
rect 8894 912 8924 946
rect 8924 912 8928 946
rect 8967 912 8992 946
rect 8992 912 9001 946
rect 9040 912 9060 946
rect 9060 912 9074 946
rect 9113 912 9128 946
rect 9128 912 9147 946
rect 9186 912 9196 946
rect 9196 912 9220 946
rect 9259 912 9264 946
rect 9264 912 9293 946
rect 9332 912 9366 946
rect 9564 912 9568 946
rect 9568 912 9598 946
rect 9637 912 9670 946
rect 9670 912 9671 946
rect 9710 912 9738 946
rect 9738 912 9744 946
rect 9783 912 9806 946
rect 9806 912 9817 946
rect 9856 912 9874 946
rect 9874 912 9890 946
rect 9929 912 9942 946
rect 9942 912 9963 946
rect 10002 912 10010 946
rect 10010 912 10036 946
rect 10075 912 10078 946
rect 10078 912 10109 946
rect 10148 912 10180 946
rect 10180 912 10182 946
rect 10221 912 10248 946
rect 10248 912 10255 946
rect 10294 912 10316 946
rect 10316 912 10328 946
rect 10367 912 10384 946
rect 10384 912 10401 946
rect 10440 912 10452 946
rect 10452 912 10474 946
rect 10514 912 10520 946
rect 10520 912 10548 946
rect 10588 912 10622 946
rect 10662 912 10690 946
rect 10690 912 10696 946
rect 10736 912 10758 946
rect 10758 912 10770 946
rect 10810 912 10826 946
rect 10826 912 10844 946
rect 10884 912 10894 946
rect 10894 912 10918 946
rect 10958 912 10962 946
rect 10962 912 10992 946
rect 11032 912 11064 946
rect 11064 912 11066 946
rect 11106 912 11132 946
rect 11132 912 11140 946
rect 11180 912 11200 946
rect 11200 912 11214 946
rect 11254 912 11268 946
rect 11268 912 11288 946
rect 11328 912 11336 946
rect 11336 912 11362 946
rect 11402 912 11404 946
rect 11404 912 11436 946
rect 11476 912 11506 946
rect 11506 912 11510 946
rect 11566 945 11599 977
rect 11599 945 11600 977
rect 7330 904 7364 905
rect 7330 871 7364 904
rect 7330 797 7364 831
rect 11566 904 11600 905
rect 11566 871 11599 904
rect 11599 871 11600 904
rect 11566 797 11599 831
rect 11599 797 11600 831
rect 7330 724 7364 757
rect 7420 756 7454 790
rect 7494 756 7496 790
rect 7496 756 7528 790
rect 7568 756 7598 790
rect 7598 756 7602 790
rect 7642 756 7666 790
rect 7666 756 7676 790
rect 7716 756 7734 790
rect 7734 756 7750 790
rect 7790 756 7802 790
rect 7802 756 7824 790
rect 7864 756 7870 790
rect 7870 756 7898 790
rect 7938 756 7972 790
rect 8012 756 8040 790
rect 8040 756 8046 790
rect 8086 756 8108 790
rect 8108 756 8120 790
rect 8160 756 8176 790
rect 8176 756 8194 790
rect 8234 756 8244 790
rect 8244 756 8268 790
rect 8308 756 8312 790
rect 8312 756 8342 790
rect 8382 756 8414 790
rect 8414 756 8416 790
rect 8456 756 8482 790
rect 8482 756 8490 790
rect 8529 756 8550 790
rect 8550 756 8563 790
rect 8602 756 8618 790
rect 8618 756 8636 790
rect 8675 756 8686 790
rect 8686 756 8709 790
rect 8748 756 8754 790
rect 8754 756 8782 790
rect 8821 756 8822 790
rect 8822 756 8855 790
rect 8894 756 8924 790
rect 8924 756 8928 790
rect 8967 756 8992 790
rect 8992 756 9001 790
rect 9040 756 9060 790
rect 9060 756 9074 790
rect 9113 756 9128 790
rect 9128 756 9147 790
rect 9186 756 9196 790
rect 9196 756 9220 790
rect 9259 756 9264 790
rect 9264 756 9293 790
rect 9332 756 9366 790
rect 9564 756 9568 790
rect 9568 756 9598 790
rect 9637 756 9670 790
rect 9670 756 9671 790
rect 9710 756 9738 790
rect 9738 756 9744 790
rect 9783 756 9806 790
rect 9806 756 9817 790
rect 9856 756 9874 790
rect 9874 756 9890 790
rect 9929 756 9942 790
rect 9942 756 9963 790
rect 10002 756 10010 790
rect 10010 756 10036 790
rect 10075 756 10078 790
rect 10078 756 10109 790
rect 10148 756 10180 790
rect 10180 756 10182 790
rect 10221 756 10248 790
rect 10248 756 10255 790
rect 10294 756 10316 790
rect 10316 756 10328 790
rect 10367 756 10384 790
rect 10384 756 10401 790
rect 10440 756 10452 790
rect 10452 756 10474 790
rect 10514 756 10520 790
rect 10520 756 10548 790
rect 10588 756 10622 790
rect 10662 756 10690 790
rect 10690 756 10696 790
rect 10736 756 10758 790
rect 10758 756 10770 790
rect 10810 756 10826 790
rect 10826 756 10844 790
rect 10884 756 10894 790
rect 10894 756 10918 790
rect 10958 756 10962 790
rect 10962 756 10992 790
rect 11032 756 11064 790
rect 11064 756 11066 790
rect 11106 756 11132 790
rect 11132 756 11140 790
rect 11180 756 11200 790
rect 11200 756 11214 790
rect 11254 756 11268 790
rect 11268 756 11288 790
rect 11328 756 11336 790
rect 11336 756 11362 790
rect 11402 756 11404 790
rect 11404 756 11436 790
rect 11476 756 11506 790
rect 11506 756 11510 790
rect 7330 723 7364 724
rect 7330 651 7364 683
rect 7330 649 7364 651
rect 11566 724 11599 757
rect 11599 724 11600 757
rect 11566 723 11600 724
rect 11566 651 11599 683
rect 11599 651 11600 683
rect 11566 649 11600 651
rect 7330 578 7364 609
rect 7420 600 7454 634
rect 7494 600 7496 634
rect 7496 600 7528 634
rect 7568 600 7598 634
rect 7598 600 7602 634
rect 7642 600 7666 634
rect 7666 600 7676 634
rect 7716 600 7734 634
rect 7734 600 7750 634
rect 7790 600 7802 634
rect 7802 600 7824 634
rect 7864 600 7870 634
rect 7870 600 7898 634
rect 7938 600 7972 634
rect 8012 600 8040 634
rect 8040 600 8046 634
rect 8086 600 8108 634
rect 8108 600 8120 634
rect 8160 600 8176 634
rect 8176 600 8194 634
rect 8234 600 8244 634
rect 8244 600 8268 634
rect 8308 600 8312 634
rect 8312 600 8342 634
rect 8382 600 8414 634
rect 8414 600 8416 634
rect 8456 600 8482 634
rect 8482 600 8490 634
rect 8529 600 8550 634
rect 8550 600 8563 634
rect 8602 600 8618 634
rect 8618 600 8636 634
rect 8675 600 8686 634
rect 8686 600 8709 634
rect 8748 600 8754 634
rect 8754 600 8782 634
rect 8821 600 8822 634
rect 8822 600 8855 634
rect 8894 600 8924 634
rect 8924 600 8928 634
rect 8967 600 8992 634
rect 8992 600 9001 634
rect 9040 600 9060 634
rect 9060 600 9074 634
rect 9113 600 9128 634
rect 9128 600 9147 634
rect 9186 600 9196 634
rect 9196 600 9220 634
rect 9259 600 9264 634
rect 9264 600 9293 634
rect 9332 600 9366 634
rect 9564 600 9568 634
rect 9568 600 9598 634
rect 9637 600 9670 634
rect 9670 600 9671 634
rect 9710 600 9738 634
rect 9738 600 9744 634
rect 9783 600 9806 634
rect 9806 600 9817 634
rect 9856 600 9874 634
rect 9874 600 9890 634
rect 9929 600 9942 634
rect 9942 600 9963 634
rect 10002 600 10010 634
rect 10010 600 10036 634
rect 10075 600 10078 634
rect 10078 600 10109 634
rect 10148 600 10180 634
rect 10180 600 10182 634
rect 10221 600 10248 634
rect 10248 600 10255 634
rect 10294 600 10316 634
rect 10316 600 10328 634
rect 10367 600 10384 634
rect 10384 600 10401 634
rect 10440 600 10452 634
rect 10452 600 10474 634
rect 10514 600 10520 634
rect 10520 600 10548 634
rect 10588 600 10622 634
rect 10662 600 10690 634
rect 10690 600 10696 634
rect 10736 600 10758 634
rect 10758 600 10770 634
rect 10810 600 10826 634
rect 10826 600 10844 634
rect 10884 600 10894 634
rect 10894 600 10918 634
rect 10958 600 10962 634
rect 10962 600 10992 634
rect 11032 600 11064 634
rect 11064 600 11066 634
rect 11106 600 11132 634
rect 11132 600 11140 634
rect 11180 600 11200 634
rect 11200 600 11214 634
rect 11254 600 11268 634
rect 11268 600 11288 634
rect 11328 600 11336 634
rect 11336 600 11362 634
rect 11402 600 11404 634
rect 11404 600 11436 634
rect 11476 600 11506 634
rect 11506 600 11510 634
rect 7330 575 7364 578
rect 7330 505 7364 535
rect 7330 501 7364 505
rect 11566 578 11599 609
rect 11599 578 11600 609
rect 11566 575 11600 578
rect 11566 505 11599 535
rect 11599 505 11600 535
rect 11566 501 11600 505
rect 11645 1312 11751 1378
rect 11645 1278 11681 1312
rect 11681 1278 11715 1312
rect 11715 1278 11751 1312
rect 11645 1244 11751 1278
rect 11645 1210 11681 1244
rect 11681 1210 11715 1244
rect 11715 1210 11751 1244
rect 11645 1200 11751 1210
rect 11645 1127 11679 1161
rect 11717 1127 11751 1161
rect 11645 1054 11679 1088
rect 11717 1054 11751 1088
rect 11645 981 11679 1015
rect 11717 981 11751 1015
rect 11645 908 11679 942
rect 11717 908 11751 942
rect 11645 835 11679 869
rect 11717 835 11751 869
rect 11645 762 11679 796
rect 11717 762 11751 796
rect 11645 689 11679 723
rect 11717 689 11751 723
rect 11645 616 11679 650
rect 11717 616 11751 650
rect 11645 543 11679 577
rect 11717 543 11751 577
rect 7420 444 7454 478
rect 7494 444 7496 478
rect 7496 444 7528 478
rect 7568 444 7598 478
rect 7598 444 7602 478
rect 7642 444 7666 478
rect 7666 444 7676 478
rect 7716 444 7734 478
rect 7734 444 7750 478
rect 7790 444 7802 478
rect 7802 444 7824 478
rect 7864 444 7870 478
rect 7870 444 7898 478
rect 7938 444 7972 478
rect 8012 444 8040 478
rect 8040 444 8046 478
rect 8086 444 8108 478
rect 8108 444 8120 478
rect 8160 444 8176 478
rect 8176 444 8194 478
rect 8234 444 8244 478
rect 8244 444 8268 478
rect 8308 444 8312 478
rect 8312 444 8342 478
rect 8382 444 8414 478
rect 8414 444 8416 478
rect 8456 444 8482 478
rect 8482 444 8490 478
rect 8529 444 8550 478
rect 8550 444 8563 478
rect 8602 444 8618 478
rect 8618 444 8636 478
rect 8675 444 8686 478
rect 8686 444 8709 478
rect 8748 444 8754 478
rect 8754 444 8782 478
rect 8821 444 8822 478
rect 8822 444 8855 478
rect 8894 444 8924 478
rect 8924 444 8928 478
rect 8967 444 8992 478
rect 8992 444 9001 478
rect 9040 444 9060 478
rect 9060 444 9074 478
rect 9113 444 9128 478
rect 9128 444 9147 478
rect 9186 444 9196 478
rect 9196 444 9220 478
rect 9259 444 9264 478
rect 9264 444 9293 478
rect 9332 444 9366 478
rect 9564 444 9568 478
rect 9568 444 9598 478
rect 9637 444 9670 478
rect 9670 444 9671 478
rect 9710 444 9738 478
rect 9738 444 9744 478
rect 9783 444 9806 478
rect 9806 444 9817 478
rect 9856 444 9874 478
rect 9874 444 9890 478
rect 9929 444 9942 478
rect 9942 444 9963 478
rect 10002 444 10010 478
rect 10010 444 10036 478
rect 10075 444 10078 478
rect 10078 444 10109 478
rect 10148 444 10180 478
rect 10180 444 10182 478
rect 10221 444 10248 478
rect 10248 444 10255 478
rect 10294 444 10316 478
rect 10316 444 10328 478
rect 10367 444 10384 478
rect 10384 444 10401 478
rect 10440 444 10452 478
rect 10452 444 10474 478
rect 10514 444 10520 478
rect 10520 444 10548 478
rect 10588 444 10622 478
rect 10662 444 10690 478
rect 10690 444 10696 478
rect 10736 444 10758 478
rect 10758 444 10770 478
rect 10810 444 10826 478
rect 10826 444 10844 478
rect 10884 444 10894 478
rect 10894 444 10918 478
rect 10958 444 10962 478
rect 10962 444 10992 478
rect 11032 444 11064 478
rect 11064 444 11066 478
rect 11106 444 11132 478
rect 11132 444 11140 478
rect 11180 444 11200 478
rect 11200 444 11214 478
rect 11254 444 11268 478
rect 11268 444 11288 478
rect 11328 444 11336 478
rect 11336 444 11362 478
rect 11402 444 11404 478
rect 11404 444 11436 478
rect 11476 444 11506 478
rect 11506 444 11510 478
rect 11645 470 11679 504
rect 11717 470 11751 504
rect 11645 397 11679 431
rect 11717 397 11751 431
rect 7163 325 7264 359
rect 7264 325 7269 359
rect 7308 325 7332 358
rect 7332 325 7342 358
rect 7381 325 7400 358
rect 7400 325 7415 358
rect 7454 325 7468 358
rect 7468 325 7488 358
rect 7527 325 7536 358
rect 7536 325 7561 358
rect 7600 325 7604 358
rect 7604 325 7634 358
rect 7673 325 7706 358
rect 7706 325 7707 358
rect 7746 325 7774 358
rect 7774 325 7780 358
rect 7819 325 7842 358
rect 7842 325 7853 358
rect 7892 325 7910 358
rect 7910 325 7926 358
rect 7965 325 7978 358
rect 7978 325 7999 358
rect 8038 325 8046 358
rect 8046 325 8072 358
rect 8111 325 8114 358
rect 8114 325 8145 358
rect 8184 325 8216 358
rect 8216 325 8218 358
rect 8257 325 8284 358
rect 8284 325 8291 358
rect 8330 325 8352 358
rect 8352 325 8364 358
rect 8403 325 8420 358
rect 8420 325 8437 358
rect 8476 325 8488 358
rect 8488 325 8510 358
rect 8549 325 8556 358
rect 8556 325 8590 358
rect 8590 325 8624 358
rect 8624 325 8658 358
rect 8658 325 8692 358
rect 8692 325 8726 358
rect 8726 325 8760 358
rect 8760 325 8794 358
rect 8794 325 8828 358
rect 8828 325 8862 358
rect 8862 325 8896 358
rect 8896 325 8930 358
rect 8930 325 8964 358
rect 8964 325 8998 358
rect 8998 325 9032 358
rect 9032 325 9066 358
rect 9066 325 9100 358
rect 9100 325 9134 358
rect 9134 325 9168 358
rect 9168 325 9202 358
rect 9202 325 9236 358
rect 9236 325 9270 358
rect 9270 325 9304 358
rect 9304 325 9338 358
rect 9338 325 9372 358
rect 9372 325 9406 358
rect 9406 325 9440 358
rect 9440 325 9474 358
rect 9474 325 9508 358
rect 9508 325 9542 358
rect 9542 325 9576 358
rect 9576 325 9610 358
rect 9610 325 9644 358
rect 9644 325 9678 358
rect 9678 325 9712 358
rect 9712 325 9746 358
rect 9746 325 9780 358
rect 9780 325 9814 358
rect 9814 325 9848 358
rect 9848 325 9882 358
rect 9882 325 9916 358
rect 9916 325 9950 358
rect 9950 325 9984 358
rect 9984 325 10018 358
rect 10018 325 10052 358
rect 10052 325 10086 358
rect 10086 325 10120 358
rect 10120 325 10154 358
rect 10154 325 10188 358
rect 10188 325 10222 358
rect 10222 325 10256 358
rect 10256 325 10290 358
rect 10290 325 10324 358
rect 10324 325 10358 358
rect 10358 325 10392 358
rect 10392 325 10426 358
rect 10426 325 10460 358
rect 10460 325 10494 358
rect 10494 325 10528 358
rect 10528 325 10562 358
rect 10562 325 10596 358
rect 10596 325 10630 358
rect 10630 325 10664 358
rect 10664 325 10698 358
rect 10698 325 10732 358
rect 10732 325 10766 358
rect 10766 325 10800 358
rect 10800 325 10834 358
rect 10834 325 10868 358
rect 10868 325 10902 358
rect 10902 325 10936 358
rect 10936 325 10970 358
rect 10970 325 11004 358
rect 11004 325 11038 358
rect 11038 325 11072 358
rect 11072 325 11106 358
rect 11106 325 11140 358
rect 11140 325 11174 358
rect 11174 325 11208 358
rect 11208 325 11242 358
rect 11242 325 11276 358
rect 11276 325 11310 358
rect 11310 325 11344 358
rect 11344 325 11378 358
rect 11378 325 11412 358
rect 11412 325 11446 358
rect 11446 325 11480 358
rect 11480 325 11514 358
rect 11514 325 11548 358
rect 11548 325 11582 358
rect 11582 325 11616 358
rect 11616 325 11650 358
rect 11650 325 11679 358
rect 7163 324 7269 325
rect 7308 324 7342 325
rect 7381 324 7415 325
rect 7454 324 7488 325
rect 7527 324 7561 325
rect 7600 324 7634 325
rect 7673 324 7707 325
rect 7746 324 7780 325
rect 7819 324 7853 325
rect 7892 324 7926 325
rect 7965 324 7999 325
rect 8038 324 8072 325
rect 8111 324 8145 325
rect 8184 324 8218 325
rect 8257 324 8291 325
rect 8330 324 8364 325
rect 8403 324 8437 325
rect 8476 324 8510 325
rect 7235 252 7269 286
rect 7308 252 7342 286
rect 7381 252 7415 286
rect 7454 252 7488 286
rect 7527 252 7561 286
rect 7600 252 7634 286
rect 7673 252 7707 286
rect 7746 252 7780 286
rect 7819 252 7853 286
rect 7892 252 7926 286
rect 7965 252 7999 286
rect 8038 252 8072 286
rect 8111 252 8145 286
rect 8184 252 8218 286
rect 8257 252 8291 286
rect 8330 252 8364 286
rect 8403 252 8437 286
rect 8476 252 8510 286
rect 8549 252 11679 325
rect 11717 324 11751 358
rect 11900 1391 11934 1425
rect 11972 1391 12006 1425
rect 11900 1318 11934 1352
rect 11972 1318 12006 1352
rect 11900 1245 11934 1279
rect 11972 1245 12006 1279
rect 11900 1172 11934 1206
rect 11972 1172 12006 1206
rect 11900 1099 11934 1133
rect 11972 1099 12006 1133
rect 11900 1025 11934 1059
rect 11972 1025 12006 1059
rect 11900 951 11934 985
rect 11972 951 12006 985
rect 11900 877 11934 911
rect 11972 877 12006 911
rect 11900 803 11934 837
rect 11972 803 12006 837
rect 11900 729 11934 763
rect 11972 729 12006 763
rect 11900 655 11934 689
rect 11972 655 12006 689
rect 11900 581 11934 615
rect 11972 581 12006 615
rect 11900 507 11934 541
rect 11972 507 12006 541
rect 11900 433 11934 467
rect 11972 433 12006 467
rect 11900 359 11934 393
rect 11972 359 12006 393
rect 11900 285 11934 319
rect 11972 285 12006 319
rect 6882 171 6988 243
rect 11900 211 11934 245
rect 11972 211 12006 245
rect 206 169 240 171
rect 279 169 313 171
rect 352 169 386 171
rect 425 169 459 171
rect 498 169 532 171
rect 571 169 605 171
rect 644 169 678 171
rect 717 169 751 171
rect 790 169 824 171
rect 863 169 897 171
rect 936 169 970 171
rect 1009 169 1043 171
rect 1082 169 1116 171
rect 1155 169 1189 171
rect 1228 169 1262 171
rect 1301 169 1335 171
rect 1374 169 1408 171
rect 1447 169 1481 171
rect 1520 169 1554 171
rect 1593 169 1627 171
rect 1666 169 1700 171
rect 1739 169 1773 171
rect 1812 169 1846 171
rect 206 137 240 169
rect 279 137 313 169
rect 352 137 386 169
rect 425 137 459 169
rect 498 137 532 169
rect 571 137 605 169
rect 644 137 678 169
rect 717 137 751 169
rect 790 137 824 169
rect 863 137 897 169
rect 936 137 970 169
rect 1009 137 1043 169
rect 1082 137 1116 169
rect 1155 137 1189 169
rect 1228 137 1262 169
rect 1301 137 1335 169
rect 1374 137 1408 169
rect 1447 137 1481 169
rect 1520 137 1554 169
rect 1593 137 1627 169
rect 1666 137 1700 169
rect 1739 137 1773 169
rect 1812 137 1846 169
rect 1885 137 1906 171
rect 1906 137 1919 171
rect 1958 137 1992 171
rect 2031 137 2065 171
rect 2104 169 2138 171
rect 2177 169 2211 171
rect 2250 169 2284 171
rect 2323 169 2357 171
rect 2396 169 11934 171
rect 2104 137 2138 169
rect 2177 137 2211 169
rect 2250 137 2284 169
rect 2323 137 2357 169
rect 133 67 138 99
rect 138 67 167 99
rect 206 67 240 99
rect 279 67 313 99
rect 352 67 386 99
rect 425 67 459 99
rect 498 67 532 99
rect 571 67 605 99
rect 644 67 678 99
rect 717 67 751 99
rect 790 67 824 99
rect 863 67 897 99
rect 936 67 970 99
rect 1009 67 1043 99
rect 1082 67 1116 99
rect 1155 67 1189 99
rect 1228 67 1262 99
rect 1301 67 1335 99
rect 1374 67 1408 99
rect 1447 67 1481 99
rect 1520 67 1554 99
rect 1593 67 1627 99
rect 1666 67 1700 99
rect 1739 67 1773 99
rect 1812 67 1846 99
rect 133 65 167 67
rect 206 65 240 67
rect 279 65 313 67
rect 352 65 386 67
rect 425 65 459 67
rect 498 65 532 67
rect 571 65 605 67
rect 644 65 678 67
rect 717 65 751 67
rect 790 65 824 67
rect 863 65 897 67
rect 936 65 970 67
rect 1009 65 1043 67
rect 1082 65 1116 67
rect 1155 65 1189 67
rect 1228 65 1262 67
rect 1301 65 1335 67
rect 1374 65 1408 67
rect 1447 65 1481 67
rect 1520 65 1554 67
rect 1593 65 1627 67
rect 1666 65 1700 67
rect 1739 65 1773 67
rect 1812 65 1846 67
rect 1885 65 1919 99
rect 1958 65 1992 99
rect 2031 67 2035 99
rect 2035 67 2065 99
rect 2104 67 2138 99
rect 2177 67 2211 99
rect 2250 67 2284 99
rect 2323 67 2357 99
rect 2396 67 4653 169
rect 4653 135 7020 169
rect 7020 135 7054 169
rect 7054 135 7089 169
rect 7089 135 7123 169
rect 7123 135 7158 169
rect 7158 135 7192 169
rect 7192 135 7227 169
rect 7227 135 7261 169
rect 7261 135 7296 169
rect 7296 135 7330 169
rect 7330 135 7365 169
rect 7365 135 7399 169
rect 7399 135 7434 169
rect 7434 135 7468 169
rect 7468 135 7503 169
rect 7503 135 7537 169
rect 7537 135 7572 169
rect 7572 135 7606 169
rect 7606 135 7641 169
rect 7641 135 7675 169
rect 7675 135 7710 169
rect 7710 135 7744 169
rect 7744 135 7779 169
rect 7779 135 7813 169
rect 7813 135 7848 169
rect 7848 135 7882 169
rect 7882 135 7917 169
rect 7917 135 7951 169
rect 7951 135 7986 169
rect 7986 135 8020 169
rect 8020 135 8055 169
rect 8055 135 8089 169
rect 8089 135 8124 169
rect 8124 135 8158 169
rect 8158 135 8193 169
rect 8193 135 8227 169
rect 8227 135 8262 169
rect 8262 135 8296 169
rect 8296 135 8331 169
rect 8331 135 8365 169
rect 8365 135 8400 169
rect 8400 135 8434 169
rect 8434 135 8469 169
rect 8469 135 8503 169
rect 8503 135 8538 169
rect 8538 135 8572 169
rect 8572 135 8607 169
rect 8607 135 8641 169
rect 8641 135 8676 169
rect 8676 135 8710 169
rect 8710 135 8745 169
rect 8745 135 8779 169
rect 8779 135 8814 169
rect 8814 135 8848 169
rect 8848 135 8883 169
rect 8883 135 8917 169
rect 8917 135 8952 169
rect 4653 101 8952 135
rect 4653 67 7020 101
rect 7020 67 7054 101
rect 7054 67 7089 101
rect 7089 67 7123 101
rect 7123 67 7158 101
rect 7158 67 7192 101
rect 7192 67 7227 101
rect 7227 67 7261 101
rect 7261 67 7296 101
rect 7296 67 7330 101
rect 7330 67 7365 101
rect 7365 67 7399 101
rect 7399 67 7434 101
rect 7434 67 7468 101
rect 7468 67 7503 101
rect 7503 67 7537 101
rect 7537 67 7572 101
rect 7572 67 7606 101
rect 7606 67 7641 101
rect 7641 67 7675 101
rect 7675 67 7710 101
rect 7710 67 7744 101
rect 7744 67 7779 101
rect 7779 67 7813 101
rect 7813 67 7848 101
rect 7848 67 7882 101
rect 7882 67 7917 101
rect 7917 67 7951 101
rect 7951 67 7986 101
rect 7986 67 8020 101
rect 8020 67 8055 101
rect 8055 67 8089 101
rect 8089 67 8124 101
rect 8124 67 8158 101
rect 8158 67 8193 101
rect 8193 67 8227 101
rect 8227 67 8262 101
rect 8262 67 8296 101
rect 8296 67 8331 101
rect 8331 67 8365 101
rect 8365 67 8400 101
rect 8400 67 8434 101
rect 8434 67 8469 101
rect 8469 67 8503 101
rect 8503 67 8538 101
rect 8538 67 8572 101
rect 8572 67 8607 101
rect 8607 67 8641 101
rect 8641 67 8676 101
rect 8676 67 8710 101
rect 8710 67 8745 101
rect 8745 67 8779 101
rect 8779 67 8814 101
rect 8814 67 8848 101
rect 8848 67 8883 101
rect 8883 67 8917 101
rect 8917 67 8952 101
rect 8952 67 11842 169
rect 11842 67 11934 169
rect 11972 137 12006 171
rect 2031 65 2065 67
rect 2104 65 2138 67
rect 2177 65 2211 67
rect 2250 65 2284 67
rect 2323 65 2357 67
rect 2396 65 11934 67
rect -496 -88 -462 -54
rect -409 -88 -375 -54
rect -322 -88 -288 -54
rect -236 -88 -202 -54
rect -150 -88 -116 -54
rect -496 -198 -462 -164
rect -409 -198 -375 -164
rect -322 -198 -288 -164
rect -236 -198 -202 -164
rect -150 -198 -116 -164
rect 5691 -1154 5725 -1153
rect 5765 -1154 5799 -1153
rect 5839 -1154 5873 -1153
rect 5913 -1154 5947 -1153
rect 5987 -1154 6021 -1153
rect 6062 -1154 6096 -1153
rect 6137 -1154 6171 -1153
rect 6212 -1154 6246 -1153
rect 6287 -1154 6321 -1153
rect 6397 -1154 6431 -1153
rect 6470 -1154 6504 -1153
rect 6543 -1154 6577 -1153
rect 5691 -1187 5698 -1154
rect 5698 -1187 5725 -1154
rect 5765 -1187 5766 -1154
rect 5766 -1187 5799 -1154
rect 5839 -1187 5868 -1154
rect 5868 -1187 5873 -1154
rect 5913 -1187 5936 -1154
rect 5936 -1187 5947 -1154
rect 5987 -1187 6004 -1154
rect 6004 -1187 6021 -1154
rect 6062 -1187 6072 -1154
rect 6072 -1187 6096 -1154
rect 6137 -1187 6140 -1154
rect 6140 -1187 6171 -1154
rect 6212 -1187 6242 -1154
rect 6242 -1187 6246 -1154
rect 6287 -1187 6310 -1154
rect 6310 -1187 6321 -1154
rect 6397 -1187 6412 -1154
rect 6412 -1187 6431 -1154
rect 6470 -1187 6480 -1154
rect 6480 -1187 6504 -1154
rect 6543 -1187 6548 -1154
rect 6548 -1187 6577 -1154
rect 6616 -1187 6650 -1153
rect 6689 -1154 6723 -1153
rect 6762 -1154 6796 -1153
rect 6835 -1154 6869 -1153
rect 6908 -1154 6942 -1153
rect 6982 -1154 7016 -1153
rect 7056 -1154 7090 -1153
rect 7130 -1154 7164 -1153
rect 7204 -1154 7238 -1153
rect 7278 -1154 7312 -1153
rect 7352 -1154 7386 -1153
rect 7426 -1154 7460 -1153
rect 6689 -1187 6718 -1154
rect 6718 -1187 6723 -1154
rect 6762 -1187 6786 -1154
rect 6786 -1187 6796 -1154
rect 6835 -1187 6854 -1154
rect 6854 -1187 6869 -1154
rect 6908 -1187 6922 -1154
rect 6922 -1187 6942 -1154
rect 6982 -1187 6990 -1154
rect 6990 -1187 7016 -1154
rect 7056 -1187 7058 -1154
rect 7058 -1187 7090 -1154
rect 7130 -1187 7160 -1154
rect 7160 -1187 7164 -1154
rect 7204 -1187 7228 -1154
rect 7228 -1187 7238 -1154
rect 7278 -1187 7296 -1154
rect 7296 -1187 7312 -1154
rect 7352 -1187 7364 -1154
rect 7364 -1187 7386 -1154
rect 7426 -1187 7432 -1154
rect 7432 -1187 7460 -1154
rect 7500 -1187 7534 -1153
rect 7574 -1154 7608 -1153
rect 7648 -1154 7682 -1153
rect 7722 -1154 7756 -1153
rect 7796 -1154 7830 -1153
rect 7870 -1154 7904 -1153
rect 7574 -1187 7602 -1154
rect 7602 -1187 7608 -1154
rect 7648 -1187 7670 -1154
rect 7670 -1187 7682 -1154
rect 7722 -1187 7738 -1154
rect 7738 -1187 7756 -1154
rect 7796 -1187 7806 -1154
rect 7806 -1187 7830 -1154
rect 7870 -1187 7874 -1154
rect 7874 -1187 7904 -1154
rect 5617 -1256 5651 -1225
rect 5617 -1259 5651 -1256
rect 5617 -1324 5651 -1304
rect 5617 -1338 5651 -1324
rect 5852 -1304 5866 -1270
rect 5866 -1304 5886 -1270
rect 5927 -1304 5934 -1270
rect 5934 -1304 5961 -1270
rect 6002 -1304 6036 -1270
rect 6077 -1304 6104 -1270
rect 6104 -1304 6111 -1270
rect 6152 -1304 6172 -1270
rect 6172 -1304 6186 -1270
rect 6227 -1304 6240 -1270
rect 6240 -1304 6261 -1270
rect 6302 -1304 6308 -1270
rect 6308 -1304 6336 -1270
rect 6377 -1304 6410 -1270
rect 6410 -1304 6411 -1270
rect 6452 -1304 6478 -1270
rect 6478 -1304 6486 -1270
rect 6527 -1304 6546 -1270
rect 6546 -1304 6561 -1270
rect 6602 -1304 6614 -1270
rect 6614 -1304 6636 -1270
rect 6676 -1304 6682 -1270
rect 6682 -1304 6710 -1270
rect 6750 -1304 6784 -1270
rect 6824 -1304 6852 -1270
rect 6852 -1304 6858 -1270
rect 6898 -1304 6920 -1270
rect 6920 -1304 6932 -1270
rect 6972 -1304 6988 -1270
rect 6988 -1304 7006 -1270
rect 7046 -1304 7056 -1270
rect 7056 -1304 7080 -1270
rect 7120 -1304 7124 -1270
rect 7124 -1304 7154 -1270
rect 7194 -1304 7226 -1270
rect 7226 -1304 7228 -1270
rect 7268 -1304 7294 -1270
rect 7294 -1304 7302 -1270
rect 7342 -1304 7362 -1270
rect 7362 -1304 7376 -1270
rect 7416 -1304 7430 -1270
rect 7430 -1304 7450 -1270
rect 7490 -1304 7498 -1270
rect 7498 -1304 7524 -1270
rect 7564 -1304 7566 -1270
rect 7566 -1304 7598 -1270
rect 7638 -1304 7668 -1270
rect 7668 -1304 7672 -1270
rect 7712 -1304 7736 -1270
rect 7736 -1304 7746 -1270
rect 7786 -1304 7804 -1270
rect 7804 -1304 7820 -1270
rect 7942 -1262 7976 -1231
rect 7942 -1265 7976 -1262
rect 5617 -1392 5651 -1383
rect 5617 -1417 5651 -1392
rect 5617 -1494 5651 -1462
rect 5617 -1496 5651 -1494
rect 5617 -1562 5651 -1541
rect 5617 -1575 5651 -1562
rect 5617 -1654 5651 -1620
rect 5617 -1724 5651 -1698
rect 5617 -1732 5651 -1724
rect 5617 -1792 5651 -1776
rect 5617 -1810 5651 -1792
rect 5617 -1860 5651 -1854
rect 5617 -1888 5651 -1860
rect 5734 -1331 5768 -1327
rect 5734 -1361 5768 -1331
rect 5734 -1402 5768 -1399
rect 5734 -1433 5768 -1402
rect 7942 -1330 7976 -1309
rect 7942 -1343 7976 -1330
rect 5852 -1460 5866 -1426
rect 5866 -1460 5886 -1426
rect 5927 -1460 5934 -1426
rect 5934 -1460 5961 -1426
rect 6002 -1460 6036 -1426
rect 6077 -1460 6104 -1426
rect 6104 -1460 6111 -1426
rect 6152 -1460 6172 -1426
rect 6172 -1460 6186 -1426
rect 6227 -1460 6240 -1426
rect 6240 -1460 6261 -1426
rect 6302 -1460 6308 -1426
rect 6308 -1460 6336 -1426
rect 6377 -1460 6410 -1426
rect 6410 -1460 6411 -1426
rect 6452 -1460 6478 -1426
rect 6478 -1460 6486 -1426
rect 6527 -1460 6546 -1426
rect 6546 -1460 6561 -1426
rect 6602 -1460 6614 -1426
rect 6614 -1460 6636 -1426
rect 6676 -1460 6682 -1426
rect 6682 -1460 6710 -1426
rect 6750 -1460 6784 -1426
rect 6824 -1460 6852 -1426
rect 6852 -1460 6858 -1426
rect 6898 -1460 6920 -1426
rect 6920 -1460 6932 -1426
rect 6972 -1460 6988 -1426
rect 6988 -1460 7006 -1426
rect 7046 -1460 7056 -1426
rect 7056 -1460 7080 -1426
rect 7120 -1460 7124 -1426
rect 7124 -1460 7154 -1426
rect 7194 -1460 7226 -1426
rect 7226 -1460 7228 -1426
rect 7268 -1460 7294 -1426
rect 7294 -1460 7302 -1426
rect 7342 -1460 7362 -1426
rect 7362 -1460 7376 -1426
rect 7416 -1460 7430 -1426
rect 7430 -1460 7450 -1426
rect 7490 -1460 7498 -1426
rect 7498 -1460 7524 -1426
rect 7564 -1460 7566 -1426
rect 7566 -1460 7598 -1426
rect 7638 -1460 7668 -1426
rect 7668 -1460 7672 -1426
rect 7712 -1460 7736 -1426
rect 7736 -1460 7746 -1426
rect 7786 -1460 7804 -1426
rect 7804 -1460 7820 -1426
rect 7942 -1398 7976 -1387
rect 7942 -1421 7976 -1398
rect 5734 -1473 5768 -1472
rect 5734 -1506 5768 -1473
rect 5734 -1579 5768 -1545
rect 7942 -1466 7976 -1465
rect 7942 -1499 7976 -1466
rect 7942 -1568 7976 -1543
rect 7942 -1577 7976 -1568
rect 5852 -1616 5866 -1582
rect 5866 -1616 5886 -1582
rect 5927 -1616 5934 -1582
rect 5934 -1616 5961 -1582
rect 6002 -1616 6036 -1582
rect 6077 -1616 6104 -1582
rect 6104 -1616 6111 -1582
rect 6152 -1616 6172 -1582
rect 6172 -1616 6186 -1582
rect 6227 -1616 6240 -1582
rect 6240 -1616 6261 -1582
rect 6302 -1616 6308 -1582
rect 6308 -1616 6336 -1582
rect 6377 -1616 6410 -1582
rect 6410 -1616 6411 -1582
rect 6452 -1616 6478 -1582
rect 6478 -1616 6486 -1582
rect 6527 -1616 6546 -1582
rect 6546 -1616 6561 -1582
rect 6602 -1616 6614 -1582
rect 6614 -1616 6636 -1582
rect 6676 -1616 6682 -1582
rect 6682 -1616 6710 -1582
rect 6750 -1616 6784 -1582
rect 6824 -1616 6852 -1582
rect 6852 -1616 6858 -1582
rect 6898 -1616 6920 -1582
rect 6920 -1616 6932 -1582
rect 6972 -1616 6988 -1582
rect 6988 -1616 7006 -1582
rect 7046 -1616 7056 -1582
rect 7056 -1616 7080 -1582
rect 7120 -1616 7124 -1582
rect 7124 -1616 7154 -1582
rect 7194 -1616 7226 -1582
rect 7226 -1616 7228 -1582
rect 7268 -1616 7294 -1582
rect 7294 -1616 7302 -1582
rect 7342 -1616 7362 -1582
rect 7362 -1616 7376 -1582
rect 7416 -1616 7430 -1582
rect 7430 -1616 7450 -1582
rect 7490 -1616 7498 -1582
rect 7498 -1616 7524 -1582
rect 7564 -1616 7566 -1582
rect 7566 -1616 7598 -1582
rect 7638 -1616 7668 -1582
rect 7668 -1616 7672 -1582
rect 7712 -1616 7736 -1582
rect 7736 -1616 7746 -1582
rect 7786 -1616 7804 -1582
rect 7804 -1616 7820 -1582
rect 5734 -1651 5768 -1618
rect 5734 -1652 5768 -1651
rect 5734 -1723 5768 -1691
rect 5734 -1725 5768 -1723
rect 7942 -1636 7976 -1622
rect 7942 -1656 7976 -1636
rect 7942 -1704 7976 -1701
rect 7942 -1735 7976 -1704
rect 5734 -1795 5768 -1764
rect 5852 -1772 5866 -1738
rect 5866 -1772 5886 -1738
rect 5927 -1772 5934 -1738
rect 5934 -1772 5961 -1738
rect 6002 -1772 6036 -1738
rect 6077 -1772 6104 -1738
rect 6104 -1772 6111 -1738
rect 6152 -1772 6172 -1738
rect 6172 -1772 6186 -1738
rect 6227 -1772 6240 -1738
rect 6240 -1772 6261 -1738
rect 6302 -1772 6308 -1738
rect 6308 -1772 6336 -1738
rect 6377 -1772 6410 -1738
rect 6410 -1772 6411 -1738
rect 6452 -1772 6478 -1738
rect 6478 -1772 6486 -1738
rect 6527 -1772 6546 -1738
rect 6546 -1772 6561 -1738
rect 6602 -1772 6614 -1738
rect 6614 -1772 6636 -1738
rect 6676 -1772 6682 -1738
rect 6682 -1772 6710 -1738
rect 6750 -1772 6784 -1738
rect 6824 -1772 6852 -1738
rect 6852 -1772 6858 -1738
rect 6898 -1772 6920 -1738
rect 6920 -1772 6932 -1738
rect 6972 -1772 6988 -1738
rect 6988 -1772 7006 -1738
rect 7046 -1772 7056 -1738
rect 7056 -1772 7080 -1738
rect 7120 -1772 7124 -1738
rect 7124 -1772 7154 -1738
rect 7194 -1772 7226 -1738
rect 7226 -1772 7228 -1738
rect 7268 -1772 7294 -1738
rect 7294 -1772 7302 -1738
rect 7342 -1772 7362 -1738
rect 7362 -1772 7376 -1738
rect 7416 -1772 7430 -1738
rect 7430 -1772 7450 -1738
rect 7490 -1772 7498 -1738
rect 7498 -1772 7524 -1738
rect 7564 -1772 7566 -1738
rect 7566 -1772 7598 -1738
rect 7638 -1772 7668 -1738
rect 7668 -1772 7672 -1738
rect 7712 -1772 7736 -1738
rect 7736 -1772 7746 -1738
rect 7786 -1772 7804 -1738
rect 7804 -1772 7820 -1738
rect 5734 -1798 5768 -1795
rect 5734 -1867 5768 -1837
rect 5734 -1871 5768 -1867
rect 7942 -1806 7976 -1780
rect 7942 -1814 7976 -1806
rect 5852 -1928 5866 -1894
rect 5866 -1928 5886 -1894
rect 5927 -1928 5934 -1894
rect 5934 -1928 5961 -1894
rect 6002 -1928 6036 -1894
rect 6077 -1928 6104 -1894
rect 6104 -1928 6111 -1894
rect 6152 -1928 6172 -1894
rect 6172 -1928 6186 -1894
rect 6227 -1928 6240 -1894
rect 6240 -1928 6261 -1894
rect 6302 -1928 6308 -1894
rect 6308 -1928 6336 -1894
rect 6377 -1928 6410 -1894
rect 6410 -1928 6411 -1894
rect 6452 -1928 6478 -1894
rect 6478 -1928 6486 -1894
rect 6527 -1928 6546 -1894
rect 6546 -1928 6561 -1894
rect 6602 -1928 6614 -1894
rect 6614 -1928 6636 -1894
rect 6676 -1928 6682 -1894
rect 6682 -1928 6710 -1894
rect 6750 -1928 6784 -1894
rect 6824 -1928 6852 -1894
rect 6852 -1928 6858 -1894
rect 6898 -1928 6920 -1894
rect 6920 -1928 6932 -1894
rect 6972 -1928 6988 -1894
rect 6988 -1928 7006 -1894
rect 7046 -1928 7056 -1894
rect 7056 -1928 7080 -1894
rect 7120 -1928 7124 -1894
rect 7124 -1928 7154 -1894
rect 7194 -1928 7226 -1894
rect 7226 -1928 7228 -1894
rect 7268 -1928 7294 -1894
rect 7294 -1928 7302 -1894
rect 7342 -1928 7362 -1894
rect 7362 -1928 7376 -1894
rect 7416 -1928 7430 -1894
rect 7430 -1928 7450 -1894
rect 7490 -1928 7498 -1894
rect 7498 -1928 7524 -1894
rect 7564 -1928 7566 -1894
rect 7566 -1928 7598 -1894
rect 7638 -1928 7668 -1894
rect 7668 -1928 7672 -1894
rect 7712 -1928 7736 -1894
rect 7736 -1928 7746 -1894
rect 7786 -1928 7804 -1894
rect 7804 -1928 7820 -1894
rect 7942 -1874 7976 -1859
rect 7942 -1893 7976 -1874
rect 5617 -1962 5651 -1932
rect 5617 -1966 5651 -1962
rect 7942 -1942 7976 -1938
rect 7942 -1972 7976 -1942
rect 5689 -2044 5719 -2010
rect 5719 -2044 5723 -2010
rect 5762 -2044 5787 -2010
rect 5787 -2044 5796 -2010
rect 5835 -2044 5855 -2010
rect 5855 -2044 5869 -2010
rect 5908 -2044 5923 -2010
rect 5923 -2044 5942 -2010
rect 5981 -2044 5991 -2010
rect 5991 -2044 6015 -2010
rect 6054 -2044 6059 -2010
rect 6059 -2044 6088 -2010
rect 6127 -2044 6161 -2010
rect 6200 -2044 6229 -2010
rect 6229 -2044 6234 -2010
rect 6273 -2044 6297 -2010
rect 6297 -2044 6307 -2010
rect 6346 -2044 6365 -2010
rect 6365 -2044 6380 -2010
rect 6419 -2044 6433 -2010
rect 6433 -2044 6453 -2010
rect 6492 -2044 6501 -2010
rect 6501 -2044 6526 -2010
rect 6565 -2044 6569 -2010
rect 6569 -2044 6599 -2010
rect 6638 -2044 6671 -2010
rect 6671 -2044 6672 -2010
rect 6711 -2044 6739 -2010
rect 6739 -2044 6745 -2010
rect 6784 -2044 6807 -2010
rect 6807 -2044 6818 -2010
rect 6857 -2044 6875 -2010
rect 6875 -2044 6891 -2010
rect 6930 -2044 6943 -2010
rect 6943 -2044 6964 -2010
rect 7003 -2044 7011 -2010
rect 7011 -2044 7037 -2010
rect 7076 -2044 7079 -2010
rect 7079 -2044 7110 -2010
rect 7149 -2044 7181 -2010
rect 7181 -2044 7183 -2010
rect 7222 -2044 7249 -2010
rect 7249 -2044 7256 -2010
rect 7294 -2044 7317 -2010
rect 7317 -2044 7328 -2010
rect 7366 -2044 7385 -2010
rect 7385 -2044 7400 -2010
rect 7438 -2044 7453 -2010
rect 7453 -2044 7472 -2010
rect 7510 -2044 7521 -2010
rect 7521 -2044 7544 -2010
rect 7582 -2044 7589 -2010
rect 7589 -2044 7616 -2010
rect 7654 -2044 7657 -2010
rect 7657 -2044 7688 -2010
rect 7726 -2044 7759 -2010
rect 7759 -2044 7760 -2010
rect 7798 -2044 7827 -2010
rect 7827 -2044 7832 -2010
rect 7870 -2044 7895 -2010
rect 7895 -2044 7904 -2010
<< metal1 >>
rect -508 1494 -104 1500
rect -508 1460 -496 1494
rect -462 1460 -409 1494
rect -375 1460 -358 1494
rect -242 1460 -236 1494
rect -202 1460 -150 1494
rect -116 1460 -104 1494
rect -508 1442 -358 1460
rect -306 1442 -294 1460
rect -242 1442 -104 1460
rect -508 1421 -104 1442
rect -508 1384 -358 1421
rect -306 1384 -294 1421
rect -242 1384 -104 1421
rect -508 1350 -496 1384
rect -462 1350 -409 1384
rect -375 1369 -358 1384
rect -242 1369 -236 1384
rect -375 1350 -322 1369
rect -288 1350 -236 1369
rect -202 1350 -150 1384
rect -116 1350 -104 1384
rect -508 1348 -104 1350
rect -508 1344 -358 1348
tri -412 1335 -403 1344 ne
rect -403 1335 -358 1344
tri -403 1301 -369 1335 ne
rect -369 1301 -358 1335
tri -369 1290 -358 1301 ne
rect -306 1296 -294 1348
rect -242 1344 -104 1348
rect 55 1408 173 1618
rect 1898 1434 2016 1618
rect 55 1374 61 1408
rect 95 1374 133 1408
rect 167 1374 173 1408
rect -242 1335 -197 1344
tri -197 1335 -188 1344 nw
rect 55 1335 173 1374
rect -242 1301 -231 1335
tri -231 1301 -197 1335 nw
rect 55 1301 61 1335
rect 95 1301 133 1335
rect 167 1301 173 1335
rect -358 1290 -242 1296
tri -242 1290 -231 1301 nw
rect 55 1262 173 1301
rect 55 1228 61 1262
rect 95 1228 133 1262
rect 167 1228 173 1262
rect 55 1189 173 1228
rect 55 1155 61 1189
rect 95 1155 133 1189
rect 167 1155 173 1189
rect 55 1116 173 1155
rect 55 1082 61 1116
rect 95 1082 133 1116
rect 167 1082 173 1116
rect -509 967 -104 1054
rect -509 851 -490 967
rect -118 851 -104 967
rect -509 792 -104 851
rect 55 1043 173 1082
rect 55 1009 61 1043
rect 95 1009 133 1043
rect 167 1009 173 1043
rect 55 970 173 1009
rect 55 936 61 970
rect 95 936 133 970
rect 167 936 173 970
rect 55 897 173 936
rect 55 863 61 897
rect 95 863 133 897
rect 167 863 173 897
rect 55 824 173 863
rect 55 790 61 824
rect 95 790 133 824
rect 167 790 173 824
rect -509 760 -104 766
rect -509 726 -497 760
rect -463 726 -410 760
rect -376 726 -323 760
rect -289 726 -236 760
rect -202 726 -150 760
rect -116 726 -104 760
rect -509 682 -104 726
rect -509 648 -497 682
rect -463 648 -410 682
rect -376 648 -323 682
rect -289 648 -236 682
rect -202 648 -150 682
rect -116 648 -104 682
rect -509 604 -104 648
rect -509 570 -497 604
rect -463 570 -410 604
rect -376 570 -323 604
rect -289 570 -236 604
rect -202 570 -150 604
rect -116 570 -104 604
rect -509 564 -104 570
rect 55 751 173 790
rect 55 717 61 751
rect 95 717 133 751
rect 167 717 173 751
rect 55 678 173 717
rect 55 644 61 678
rect 95 644 133 678
rect 167 644 173 678
rect 55 605 173 644
rect 55 571 61 605
rect 95 571 133 605
rect 167 571 173 605
rect 55 532 173 571
rect 55 498 61 532
rect 95 498 133 532
rect 167 498 173 532
rect 55 459 173 498
rect 55 137 61 459
rect 167 209 173 459
rect 318 1426 1748 1432
rect 318 1392 402 1426
rect 436 1392 480 1426
rect 514 1392 558 1426
rect 592 1392 636 1426
rect 670 1392 714 1426
rect 748 1392 792 1426
rect 826 1392 870 1426
rect 904 1392 949 1426
rect 983 1392 1059 1426
rect 318 1354 1059 1392
rect 318 1320 324 1354
rect 358 1320 396 1354
rect 430 1320 480 1354
rect 514 1320 558 1354
rect 592 1320 636 1354
rect 670 1320 714 1354
rect 748 1320 792 1354
rect 826 1320 870 1354
rect 904 1320 949 1354
rect 983 1320 1059 1354
rect 1597 1392 1636 1426
rect 1670 1392 1748 1426
rect 1597 1354 1748 1392
rect 1597 1320 1636 1354
rect 1670 1350 1748 1354
rect 1670 1320 1708 1350
rect 318 1316 1708 1320
rect 1742 1316 1748 1350
rect 318 1314 1748 1316
rect 318 1305 467 1314
tri 467 1305 476 1314 nw
tri 1590 1305 1599 1314 ne
rect 1599 1305 1748 1314
rect 318 1284 446 1305
tri 446 1284 467 1305 nw
tri 1599 1284 1620 1305 ne
rect 1620 1284 1748 1305
rect 318 1277 436 1284
rect 318 1243 324 1277
rect 358 1243 396 1277
rect 430 1243 436 1277
tri 436 1274 446 1284 nw
tri 1620 1274 1630 1284 ne
rect 1630 1274 1748 1284
rect 318 1200 436 1243
rect 318 1166 324 1200
rect 358 1166 396 1200
rect 430 1166 436 1200
rect 554 1235 1504 1241
rect 554 1201 566 1235
rect 600 1201 641 1235
rect 675 1201 716 1235
rect 750 1201 791 1235
rect 825 1201 866 1235
rect 900 1201 940 1235
rect 974 1201 1014 1235
rect 1048 1201 1088 1235
rect 1122 1201 1162 1235
rect 1196 1201 1236 1235
rect 1270 1201 1310 1235
rect 1344 1201 1384 1235
rect 1418 1201 1458 1235
rect 1492 1201 1504 1235
rect 554 1195 1504 1201
rect 1630 1240 1636 1274
rect 1670 1240 1708 1274
rect 1742 1240 1748 1274
rect 1630 1198 1748 1240
tri 606 1187 614 1195 ne
rect 614 1187 933 1195
tri 933 1187 941 1195 nw
rect 318 1123 436 1166
rect 318 1089 324 1123
rect 358 1089 396 1123
rect 430 1089 436 1123
rect 318 1046 436 1089
rect 318 1012 324 1046
rect 358 1012 396 1046
rect 430 1012 436 1046
rect 318 969 436 1012
rect 318 967 324 969
rect 358 967 396 969
rect 430 967 436 969
rect 318 851 320 967
rect 318 816 436 851
rect 318 782 324 816
rect 358 782 396 816
rect 430 782 436 816
rect 318 740 436 782
rect 318 706 324 740
rect 358 706 396 740
rect 430 706 436 740
rect 318 664 436 706
rect 318 630 324 664
rect 358 630 396 664
rect 430 630 436 664
rect 318 588 436 630
rect 318 554 324 588
rect 358 554 396 588
rect 430 554 436 588
rect 318 512 436 554
rect 318 478 324 512
rect 358 478 396 512
rect 430 478 436 512
rect 318 436 436 478
rect 467 1175 519 1187
rect 467 1141 476 1175
rect 510 1141 519 1175
tri 614 1167 634 1187 ne
rect 467 1102 519 1141
rect 467 1068 476 1102
rect 510 1068 519 1102
rect 467 1029 519 1068
rect 467 995 476 1029
rect 510 995 519 1029
rect 467 956 519 995
rect 467 922 476 956
rect 510 922 519 956
rect 634 1143 913 1187
tri 913 1167 933 1187 nw
rect 634 1091 640 1143
rect 692 1091 712 1143
rect 764 1091 784 1143
rect 836 1091 855 1143
rect 907 1091 913 1143
rect 1630 1164 1636 1198
rect 1670 1164 1708 1198
rect 1742 1164 1748 1198
rect 634 1079 913 1091
rect 634 1027 640 1079
rect 692 1027 712 1079
rect 764 1027 784 1079
rect 836 1027 855 1079
rect 907 1027 913 1079
tri 615 936 634 955 se
rect 634 936 913 1027
rect 1112 1081 1118 1133
rect 1170 1081 1195 1133
rect 1247 1081 1272 1133
rect 1324 1081 1348 1133
rect 1400 1081 1424 1133
rect 1476 1081 1500 1133
rect 1552 1081 1558 1133
rect 1112 1076 1558 1081
rect 1112 1055 1124 1076
rect 1158 1055 1202 1076
rect 1236 1055 1280 1076
rect 1314 1055 1358 1076
rect 1392 1055 1435 1076
rect 1469 1055 1512 1076
rect 1546 1055 1558 1076
rect 1112 1003 1118 1055
rect 1170 1003 1195 1055
rect 1247 1003 1272 1055
rect 1324 1003 1348 1055
rect 1400 1003 1424 1055
rect 1476 1003 1500 1055
rect 1552 1003 1558 1055
rect 1630 1122 1748 1164
rect 1630 1088 1636 1122
rect 1670 1088 1708 1122
rect 1742 1088 1748 1122
rect 1630 1046 1748 1088
rect 1630 1012 1636 1046
rect 1670 1012 1708 1046
rect 1742 1012 1748 1046
rect 1630 970 1748 1012
tri 913 936 933 956 sw
rect 1630 936 1636 970
rect 1670 936 1708 970
rect 1742 936 1748 970
tri 606 927 615 936 se
rect 615 927 933 936
tri 933 927 942 936 sw
rect 467 883 519 922
rect 467 849 476 883
rect 510 849 519 883
rect 554 921 1504 927
rect 554 887 566 921
rect 600 887 641 921
rect 675 887 716 921
rect 750 887 791 921
rect 825 887 866 921
rect 900 887 940 921
rect 974 887 1014 921
rect 1048 887 1088 921
rect 1122 887 1162 921
rect 1196 887 1236 921
rect 1270 887 1310 921
rect 1344 887 1384 921
rect 1418 887 1458 921
rect 1492 887 1504 921
rect 554 881 1504 887
rect 1630 894 1748 936
rect 467 810 519 849
rect 467 776 476 810
rect 510 776 519 810
rect 1630 860 1636 894
rect 1670 860 1708 894
rect 1742 860 1748 894
rect 1630 818 1748 860
rect 467 738 519 776
rect 554 790 640 796
rect 554 756 566 790
rect 600 756 640 790
rect 554 750 640 756
tri 591 741 600 750 ne
rect 600 744 640 750
rect 692 744 712 796
rect 764 744 784 796
rect 836 744 855 796
rect 907 790 1504 796
rect 907 756 940 790
rect 974 756 1014 790
rect 1048 756 1088 790
rect 1122 756 1162 790
rect 1196 756 1236 790
rect 1270 756 1310 790
rect 1344 756 1384 790
rect 1418 756 1458 790
rect 1492 756 1504 790
rect 907 750 1504 756
rect 1630 784 1636 818
rect 1670 784 1708 818
rect 1742 784 1748 818
rect 907 744 933 750
rect 600 741 933 744
tri 933 741 942 750 nw
rect 1630 741 1748 784
rect 467 704 476 738
rect 510 704 519 738
tri 600 722 619 741 ne
rect 619 732 914 741
rect 619 722 640 732
tri 619 712 629 722 ne
rect 467 666 519 704
rect 467 632 476 666
rect 510 632 519 666
rect 467 598 519 632
rect 467 534 519 546
rect 629 680 640 722
rect 692 680 712 732
rect 764 680 784 732
rect 836 680 855 732
rect 907 680 914 732
tri 914 722 933 741 nw
rect 1630 707 1636 741
rect 1670 707 1708 741
rect 1742 707 1748 741
tri 627 510 629 512 se
rect 629 510 914 680
rect 1111 630 1117 682
rect 1169 630 1194 682
rect 1246 630 1271 682
rect 1323 630 1348 682
rect 1400 630 1424 682
rect 1476 630 1500 682
rect 1552 630 1558 682
rect 1111 604 1123 630
rect 1157 604 1201 630
rect 1235 604 1279 630
rect 1313 604 1357 630
rect 1391 604 1435 630
rect 1469 604 1512 630
rect 1546 604 1558 630
rect 1111 552 1117 604
rect 1169 552 1194 604
rect 1246 552 1271 604
rect 1323 552 1348 604
rect 1400 552 1424 604
rect 1476 552 1500 604
rect 1552 552 1558 604
rect 1630 664 1748 707
rect 1630 630 1636 664
rect 1670 630 1708 664
rect 1742 630 1748 664
rect 1630 587 1748 630
rect 1630 553 1636 587
rect 1670 553 1708 587
rect 1742 553 1748 587
tri 914 510 916 512 sw
rect 1630 510 1748 553
tri 601 484 627 510 se
rect 627 484 916 510
tri 916 484 942 510 sw
rect 467 476 519 482
rect 554 478 1504 484
rect 554 444 566 478
rect 600 444 641 478
rect 675 444 716 478
rect 750 444 791 478
rect 825 444 866 478
rect 900 444 940 478
rect 974 444 1014 478
rect 1048 444 1088 478
rect 1122 444 1162 478
rect 1196 444 1236 478
rect 1270 444 1310 478
rect 1344 444 1384 478
rect 1418 444 1458 478
rect 1492 444 1504 478
rect 554 438 1504 444
rect 1630 476 1636 510
rect 1670 476 1708 510
rect 1742 476 1748 510
rect 318 402 324 436
rect 358 402 396 436
rect 430 402 436 436
rect 1630 433 1748 476
rect 318 399 436 402
tri 436 399 439 402 sw
tri 1627 399 1630 402 se
rect 1630 399 1636 433
rect 1670 399 1708 433
rect 1742 399 1748 433
rect 318 391 439 399
tri 439 391 447 399 sw
tri 1619 391 1627 399 se
rect 1627 391 1748 399
rect 318 362 447 391
tri 447 362 476 391 sw
tri 1590 362 1619 391 se
rect 1619 362 1748 391
rect 318 360 1748 362
rect 318 326 324 360
rect 358 356 1748 360
rect 358 326 396 356
rect 318 322 396 326
rect 430 322 469 356
rect 503 322 542 356
rect 576 322 615 356
rect 649 322 688 356
rect 722 322 761 356
rect 795 322 834 356
rect 868 322 907 356
rect 941 322 980 356
rect 1014 322 1053 356
rect 1087 322 1126 356
rect 1160 322 1199 356
rect 1233 322 1272 356
rect 1306 322 1345 356
rect 1379 322 1418 356
rect 1452 322 1491 356
rect 1525 322 1564 356
rect 318 284 1564 322
rect 318 250 396 284
rect 430 250 469 284
rect 503 250 542 284
rect 576 250 615 284
rect 649 250 688 284
rect 722 250 761 284
rect 795 250 834 284
rect 868 250 907 284
rect 941 250 980 284
rect 1014 250 1053 284
rect 1087 250 1126 284
rect 1160 250 1199 284
rect 1233 250 1272 284
rect 1306 250 1345 284
rect 1379 250 1418 284
rect 1452 250 1491 284
rect 1525 250 1564 284
rect 1670 322 1708 356
rect 1742 322 1748 356
rect 1670 250 1748 322
rect 318 244 1748 250
rect 1898 1400 1904 1434
rect 1938 1400 1976 1434
rect 2010 1400 2016 1434
rect 1898 1359 2016 1400
rect 1898 1325 1904 1359
rect 1938 1325 1976 1359
rect 2010 1325 2016 1359
rect 1898 1284 2016 1325
rect 1898 1250 1904 1284
rect 1938 1250 1976 1284
rect 2010 1250 2016 1284
rect 1898 1209 2016 1250
rect 1898 1175 1904 1209
rect 1938 1175 1976 1209
rect 2010 1175 2016 1209
rect 1898 1134 2016 1175
rect 1898 1100 1904 1134
rect 1938 1100 1976 1134
rect 2010 1100 2016 1134
rect 1898 1059 2016 1100
rect 1898 1025 1904 1059
rect 1938 1025 1976 1059
rect 2010 1025 2016 1059
rect 1898 984 2016 1025
rect 1898 950 1904 984
rect 1938 950 1976 984
rect 2010 950 2016 984
rect 1898 909 2016 950
rect 1898 875 1904 909
rect 1938 875 1976 909
rect 2010 875 2016 909
rect 1898 835 2016 875
rect 1898 801 1904 835
rect 1938 801 1976 835
rect 2010 801 2016 835
rect 1898 761 2016 801
rect 1898 727 1904 761
rect 1938 727 1976 761
rect 2010 727 2016 761
rect 1898 687 2016 727
rect 1898 653 1904 687
rect 1938 653 1976 687
rect 2010 653 2016 687
rect 1898 613 2016 653
rect 1898 579 1904 613
rect 1938 579 1976 613
rect 2010 579 2016 613
rect 1898 539 2016 579
rect 1898 505 1904 539
rect 1938 505 1976 539
rect 2010 505 2016 539
rect 1898 465 2016 505
rect 1898 431 1904 465
rect 1938 431 1976 465
rect 2010 431 2016 465
rect 1898 391 2016 431
rect 1898 357 1904 391
rect 1938 357 1976 391
rect 2010 357 2016 391
rect 1898 317 2016 357
rect 1898 283 1904 317
rect 1938 283 1976 317
rect 2010 283 2016 317
rect 1898 243 2016 283
rect 2153 1450 3599 1456
rect 3651 1450 3665 1456
rect 3717 1450 3731 1456
rect 3783 1450 3797 1456
rect 3849 1450 3863 1456
rect 3915 1450 3929 1456
rect 3981 1450 3995 1456
rect 2153 1416 2237 1450
rect 2271 1416 2315 1450
rect 2349 1416 2393 1450
rect 2427 1416 2471 1450
rect 2505 1416 2549 1450
rect 2583 1416 2627 1450
rect 2661 1416 2705 1450
rect 2739 1416 2784 1450
rect 2818 1416 2894 1450
rect 2928 1416 2967 1450
rect 3001 1416 3040 1450
rect 3074 1416 3113 1450
rect 3147 1416 3186 1450
rect 3220 1416 3259 1450
rect 3293 1416 3332 1450
rect 3366 1416 3405 1450
rect 3439 1416 3478 1450
rect 3512 1416 3551 1450
rect 3585 1416 3599 1450
rect 3658 1416 3665 1450
rect 3915 1416 3916 1450
rect 3981 1416 3989 1450
rect 2153 1404 3599 1416
rect 3651 1404 3665 1416
rect 3717 1404 3731 1416
rect 3783 1404 3797 1416
rect 3849 1404 3863 1416
rect 3915 1404 3929 1416
rect 3981 1404 3995 1416
rect 4047 1404 4061 1456
rect 4113 1404 4127 1456
rect 4179 1404 4193 1456
rect 4245 1404 4259 1456
rect 4311 1450 4325 1456
rect 4377 1450 4391 1456
rect 4443 1450 4457 1456
rect 4509 1450 4523 1456
rect 4575 1450 4589 1456
rect 4641 1450 4655 1456
rect 4707 1450 4721 1456
rect 4315 1416 4325 1450
rect 4388 1416 4391 1450
rect 4641 1416 4646 1450
rect 4707 1416 4719 1450
rect 4311 1404 4325 1416
rect 4377 1404 4391 1416
rect 4443 1404 4457 1416
rect 4509 1404 4523 1416
rect 4575 1404 4589 1416
rect 4641 1404 4655 1416
rect 4707 1404 4721 1416
rect 4773 1404 4786 1456
rect 4838 1404 4851 1456
rect 4903 1404 4916 1456
rect 4968 1450 4981 1456
rect 5033 1450 5046 1456
rect 5098 1450 5111 1456
rect 5163 1450 5176 1456
rect 5228 1450 5241 1456
rect 5293 1450 6840 1456
rect 4972 1416 4981 1450
rect 5045 1416 5046 1450
rect 5228 1416 5230 1450
rect 5293 1416 5303 1450
rect 5337 1416 5376 1450
rect 5410 1416 5449 1450
rect 5483 1416 5522 1450
rect 5556 1416 5595 1450
rect 5629 1416 5668 1450
rect 5702 1416 5741 1450
rect 5775 1416 5814 1450
rect 5848 1416 5887 1450
rect 5921 1416 5961 1450
rect 5995 1416 6035 1450
rect 6069 1416 6109 1450
rect 6143 1416 6183 1450
rect 6217 1416 6257 1450
rect 6291 1416 6331 1450
rect 6365 1416 6405 1450
rect 6439 1416 6479 1450
rect 6513 1416 6553 1450
rect 6587 1416 6627 1450
rect 4968 1404 4981 1416
rect 5033 1404 5046 1416
rect 5098 1404 5111 1416
rect 5163 1404 5176 1416
rect 5228 1404 5241 1416
rect 5293 1404 6644 1416
rect 2153 1398 6644 1404
rect 6696 1398 6716 1450
rect 6768 1398 6788 1450
rect 2153 1392 6840 1398
rect 2153 1378 3599 1392
rect 3651 1378 3665 1392
rect 3717 1378 3731 1392
rect 3783 1378 3797 1392
rect 3849 1378 3863 1392
rect 3915 1378 3929 1392
rect 3981 1378 3995 1392
rect 2153 1344 2159 1378
rect 2193 1344 2231 1378
rect 2265 1344 2315 1378
rect 2349 1344 2393 1378
rect 2427 1344 2471 1378
rect 2505 1344 2549 1378
rect 2583 1344 2627 1378
rect 2661 1344 2705 1378
rect 2739 1344 2784 1378
rect 2818 1344 2894 1378
rect 2928 1344 2967 1378
rect 3001 1344 3040 1378
rect 3074 1344 3113 1378
rect 3147 1344 3186 1378
rect 3220 1344 3259 1378
rect 3293 1344 3332 1378
rect 3366 1344 3405 1378
rect 3439 1344 3478 1378
rect 3512 1344 3551 1378
rect 3585 1344 3599 1378
rect 3658 1344 3665 1378
rect 3915 1344 3916 1378
rect 3981 1344 3989 1378
rect 2153 1340 3599 1344
rect 3651 1340 3665 1344
rect 3717 1340 3731 1344
rect 3783 1340 3797 1344
rect 3849 1340 3863 1344
rect 3915 1340 3929 1344
rect 3981 1340 3995 1344
rect 4047 1340 4061 1392
rect 4113 1340 4127 1392
rect 4179 1340 4193 1392
rect 4245 1340 4259 1392
rect 4311 1378 4325 1392
rect 4377 1378 4391 1392
rect 4443 1378 4457 1392
rect 4509 1378 4523 1392
rect 4575 1378 4589 1392
rect 4641 1378 4655 1392
rect 4707 1378 4721 1392
rect 4315 1344 4325 1378
rect 4388 1344 4391 1378
rect 4641 1344 4646 1378
rect 4707 1344 4719 1378
rect 4311 1340 4325 1344
rect 4377 1340 4391 1344
rect 4443 1340 4457 1344
rect 4509 1340 4523 1344
rect 4575 1340 4589 1344
rect 4641 1340 4655 1344
rect 4707 1340 4721 1344
rect 4773 1340 4786 1392
rect 4838 1340 4851 1392
rect 4903 1340 4916 1392
rect 4968 1378 4981 1392
rect 5033 1378 5046 1392
rect 5098 1378 5111 1392
rect 5163 1378 5176 1392
rect 5228 1378 5241 1392
rect 5293 1379 6840 1392
rect 5293 1378 6644 1379
rect 6696 1378 6716 1379
rect 4972 1344 4981 1378
rect 5045 1344 5046 1378
rect 5228 1344 5230 1378
rect 5293 1344 5303 1378
rect 5337 1344 5376 1378
rect 5410 1344 5449 1378
rect 5483 1344 5522 1378
rect 5556 1344 5595 1378
rect 5629 1344 5668 1378
rect 5702 1344 5741 1378
rect 5775 1344 5814 1378
rect 5848 1344 5887 1378
rect 5921 1344 5961 1378
rect 5995 1344 6035 1378
rect 6069 1344 6109 1378
rect 6143 1344 6183 1378
rect 6217 1344 6257 1378
rect 6291 1344 6331 1378
rect 6365 1344 6405 1378
rect 6439 1344 6479 1378
rect 6513 1344 6553 1378
rect 6587 1344 6627 1378
rect 4968 1340 4981 1344
rect 5033 1340 5046 1344
rect 5098 1340 5111 1344
rect 5163 1340 5176 1344
rect 5228 1340 5241 1344
rect 5293 1340 6627 1344
rect 2153 1338 6627 1340
rect 2153 1321 2294 1338
tri 2294 1321 2311 1338 nw
tri 6566 1321 6583 1338 ne
rect 6583 1321 6627 1338
rect 6768 1327 6788 1379
rect 2153 1305 2271 1321
rect 2153 1271 2159 1305
rect 2193 1271 2231 1305
rect 2265 1271 2271 1305
tri 2271 1298 2294 1321 nw
tri 6583 1298 6606 1321 ne
rect 6606 1298 6627 1321
tri 6606 1283 6621 1298 ne
rect 2153 1232 2271 1271
tri 3127 1264 3130 1267 se
rect 3130 1264 3136 1267
rect 2153 1198 2159 1232
rect 2193 1198 2231 1232
rect 2265 1198 2271 1232
rect 2389 1258 3136 1264
rect 2389 1224 2401 1258
rect 2435 1224 2475 1258
rect 2509 1224 2549 1258
rect 2583 1224 2623 1258
rect 2657 1224 2697 1258
rect 2731 1224 2771 1258
rect 2805 1224 2845 1258
rect 2879 1224 2919 1258
rect 2953 1224 2993 1258
rect 3027 1224 3067 1258
rect 3101 1224 3136 1258
rect 2389 1218 3136 1224
tri 3127 1215 3130 1218 ne
rect 3130 1215 3136 1218
rect 3188 1215 3203 1267
rect 3255 1215 3269 1267
rect 3321 1258 3335 1267
rect 3387 1258 3401 1267
rect 3453 1264 3459 1267
tri 3459 1264 3462 1267 sw
rect 3453 1258 4359 1264
rect 3323 1224 3335 1258
rect 3397 1224 3401 1258
rect 3471 1224 3510 1258
rect 3544 1224 3583 1258
rect 3617 1224 3656 1258
rect 3690 1224 3729 1258
rect 3763 1224 3802 1258
rect 3836 1224 3875 1258
rect 3909 1224 3948 1258
rect 3982 1224 4021 1258
rect 4055 1224 4094 1258
rect 4128 1224 4167 1258
rect 4201 1224 4240 1258
rect 4274 1224 4313 1258
rect 4347 1224 4359 1258
rect 3321 1215 3335 1224
rect 3387 1215 3401 1224
rect 3453 1218 4359 1224
rect 4533 1258 5820 1267
rect 5872 1258 5885 1267
rect 5937 1258 5949 1267
rect 4533 1224 4545 1258
rect 4579 1224 4618 1258
rect 4652 1224 4691 1258
rect 4725 1224 4764 1258
rect 4798 1224 4837 1258
rect 4871 1224 4910 1258
rect 4944 1224 4983 1258
rect 5017 1224 5056 1258
rect 5090 1224 5129 1258
rect 5163 1224 5202 1258
rect 5236 1224 5275 1258
rect 5309 1224 5348 1258
rect 5382 1224 5421 1258
rect 5455 1224 5495 1258
rect 5529 1224 5569 1258
rect 5603 1224 5643 1258
rect 5677 1224 5717 1258
rect 5751 1224 5791 1258
rect 5937 1224 5939 1258
rect 3453 1215 3459 1218
tri 3459 1215 3462 1218 nw
rect 4533 1215 5820 1224
rect 5872 1215 5885 1224
rect 5937 1215 5949 1224
rect 6001 1215 6013 1267
rect 6065 1215 6077 1267
rect 6129 1215 6141 1267
rect 6193 1258 6205 1267
rect 6257 1258 6269 1267
rect 6321 1258 6333 1267
rect 6385 1258 6397 1267
rect 6449 1258 6503 1267
rect 6195 1224 6205 1258
rect 6449 1224 6457 1258
rect 6491 1224 6503 1258
rect 6193 1215 6205 1224
rect 6257 1215 6269 1224
rect 6321 1215 6333 1224
rect 6385 1215 6397 1224
rect 6449 1215 6503 1224
rect 6539 1264 6591 1270
rect 2153 1159 2271 1198
rect 2153 1141 2159 1159
rect 2193 1141 2231 1159
rect 2265 1141 2271 1159
rect 2153 1089 2154 1141
rect 2206 1089 2218 1141
rect 2270 1089 2271 1141
rect 2153 1086 2271 1089
rect 2153 1075 2159 1086
rect 2193 1075 2231 1086
rect 2265 1075 2271 1086
rect 2153 1023 2154 1075
rect 2206 1023 2218 1075
rect 2270 1023 2271 1075
rect 2153 1013 2271 1023
rect 2153 1009 2159 1013
rect 2193 1009 2231 1013
rect 2265 1009 2271 1013
rect 2153 957 2154 1009
rect 2206 957 2218 1009
rect 2270 957 2271 1009
rect 2153 940 2271 957
rect 2153 906 2159 940
rect 2193 906 2231 940
rect 2265 906 2271 940
rect 2153 867 2271 906
rect 2153 833 2159 867
rect 2193 833 2231 867
rect 2265 833 2271 867
rect 2153 794 2271 833
rect 2153 760 2159 794
rect 2193 760 2231 794
rect 2265 760 2271 794
rect 2153 721 2271 760
rect 2153 687 2159 721
rect 2193 687 2231 721
rect 2265 687 2271 721
rect 2153 648 2271 687
rect 2153 614 2159 648
rect 2193 614 2231 648
rect 2265 614 2271 648
rect 2305 1207 2357 1213
rect 2305 1134 2357 1155
rect 6539 1201 6591 1212
rect 6539 1191 6547 1201
rect 6581 1191 6591 1201
rect 6539 1133 6591 1139
rect 6621 1200 6627 1298
rect 6733 1200 6840 1327
rect 6621 1161 6840 1200
rect 6541 1129 6587 1133
tri 3590 1108 3593 1111 se
rect 3593 1108 3599 1111
rect 2305 1061 2357 1082
rect 2389 1102 3599 1108
rect 3651 1102 3670 1111
rect 3722 1102 3741 1111
rect 3793 1102 3811 1111
rect 3863 1102 3881 1111
rect 3933 1102 3951 1111
rect 2389 1068 2401 1102
rect 2435 1068 2475 1102
rect 2509 1068 2549 1102
rect 2583 1068 2623 1102
rect 2657 1068 2697 1102
rect 2731 1068 2771 1102
rect 2805 1068 2845 1102
rect 2879 1068 2919 1102
rect 2953 1068 2993 1102
rect 3027 1068 3067 1102
rect 3101 1068 3141 1102
rect 3175 1068 3215 1102
rect 3249 1068 3289 1102
rect 3323 1068 3363 1102
rect 3397 1068 3437 1102
rect 3471 1068 3510 1102
rect 3544 1068 3583 1102
rect 3651 1068 3656 1102
rect 3722 1068 3729 1102
rect 3793 1068 3802 1102
rect 3863 1068 3875 1102
rect 3933 1068 3948 1102
rect 2389 1062 3599 1068
tri 3590 1059 3593 1062 ne
rect 3593 1059 3599 1062
rect 3651 1059 3670 1068
rect 3722 1059 3741 1068
rect 3793 1059 3811 1068
rect 3863 1059 3881 1068
rect 3933 1059 3951 1068
rect 4003 1059 4021 1111
rect 4073 1059 4091 1111
rect 4143 1059 4161 1111
rect 4213 1059 4231 1111
rect 4283 1059 4301 1111
rect 4353 1059 4359 1111
rect 4533 1059 4539 1111
rect 4591 1059 4609 1111
rect 4661 1059 4679 1111
rect 4731 1059 4749 1111
rect 4801 1059 4819 1111
rect 4871 1059 4889 1111
rect 4941 1102 4959 1111
rect 5011 1102 5029 1111
rect 5081 1102 5099 1111
rect 5151 1102 5170 1111
rect 5222 1102 5241 1111
rect 5293 1102 6162 1111
rect 6214 1102 6250 1111
rect 6302 1102 6338 1111
rect 6390 1102 6503 1111
rect 4944 1068 4959 1102
rect 5017 1068 5029 1102
rect 5090 1068 5099 1102
rect 5163 1068 5170 1102
rect 5236 1068 5241 1102
rect 5309 1068 5348 1102
rect 5382 1068 5421 1102
rect 5455 1068 5495 1102
rect 5529 1068 5569 1102
rect 5603 1068 5643 1102
rect 5677 1068 5717 1102
rect 5751 1068 5791 1102
rect 5825 1068 5865 1102
rect 5899 1068 5939 1102
rect 5973 1068 6013 1102
rect 6047 1068 6087 1102
rect 6121 1068 6161 1102
rect 6214 1068 6235 1102
rect 6302 1068 6309 1102
rect 6417 1068 6457 1102
rect 6491 1068 6503 1102
rect 4941 1059 4959 1068
rect 5011 1059 5029 1068
rect 5081 1059 5099 1068
rect 5151 1059 5170 1068
rect 5222 1059 5241 1068
rect 5293 1059 6162 1068
rect 6214 1059 6250 1068
rect 6302 1059 6338 1068
rect 6390 1059 6503 1068
rect 6541 1095 6547 1129
rect 6581 1095 6587 1129
rect 2305 988 2357 1009
rect 6541 1056 6587 1095
rect 6541 1022 6547 1056
rect 6581 1022 6587 1056
rect 6541 983 6587 1022
tri 3127 952 3130 955 se
rect 3130 952 3136 955
rect 2305 915 2357 936
rect 2389 946 3136 952
rect 2389 912 2401 946
rect 2435 912 2475 946
rect 2509 912 2549 946
rect 2583 912 2623 946
rect 2657 912 2697 946
rect 2731 912 2771 946
rect 2805 912 2845 946
rect 2879 912 2919 946
rect 2953 912 2993 946
rect 3027 912 3067 946
rect 3101 912 3136 946
rect 2389 906 3136 912
tri 3127 903 3130 906 ne
rect 3130 903 3136 906
rect 3188 903 3203 955
rect 3255 903 3269 955
rect 3321 946 3335 955
rect 3387 946 3401 955
rect 3453 952 3459 955
tri 3459 952 3462 955 sw
rect 3453 946 4359 952
rect 3323 912 3335 946
rect 3397 912 3401 946
rect 3471 912 3510 946
rect 3544 912 3583 946
rect 3617 912 3656 946
rect 3690 912 3729 946
rect 3763 912 3802 946
rect 3836 912 3875 946
rect 3909 912 3948 946
rect 3982 912 4021 946
rect 4055 912 4094 946
rect 4128 912 4167 946
rect 4201 912 4240 946
rect 4274 912 4313 946
rect 4347 912 4359 946
rect 3321 903 3335 912
rect 3387 903 3401 912
rect 3453 906 4359 912
rect 4533 946 5820 955
rect 5872 946 5885 955
rect 5937 946 5949 955
rect 4533 912 4545 946
rect 4579 912 4618 946
rect 4652 912 4691 946
rect 4725 912 4764 946
rect 4798 912 4837 946
rect 4871 912 4910 946
rect 4944 912 4983 946
rect 5017 912 5056 946
rect 5090 912 5129 946
rect 5163 912 5202 946
rect 5236 912 5275 946
rect 5309 912 5348 946
rect 5382 912 5421 946
rect 5455 912 5495 946
rect 5529 912 5569 946
rect 5603 912 5643 946
rect 5677 912 5717 946
rect 5751 912 5791 946
rect 5937 912 5939 946
rect 3453 903 3459 906
tri 3459 903 3462 906 nw
rect 4533 903 5820 912
rect 5872 903 5885 912
rect 5937 903 5949 912
rect 6001 903 6013 955
rect 6065 903 6077 955
rect 6129 903 6141 955
rect 6193 946 6205 955
rect 6257 946 6269 955
rect 6321 946 6333 955
rect 6385 946 6397 955
rect 6449 946 6503 955
rect 6195 912 6205 946
rect 6449 912 6457 946
rect 6491 912 6503 946
rect 6193 903 6205 912
rect 6257 903 6269 912
rect 6321 903 6333 912
rect 6385 903 6397 912
rect 6449 903 6503 912
rect 6541 949 6547 983
rect 6581 949 6587 983
rect 6541 910 6587 949
rect 2305 842 2357 863
rect 6541 876 6547 910
rect 6581 876 6587 910
rect 6541 837 6587 876
rect 6541 803 6547 837
rect 6581 803 6587 837
tri 3592 798 3593 799 se
rect 3593 798 3599 799
tri 3591 797 3592 798 se
rect 3592 797 3599 798
tri 3590 796 3591 797 se
rect 3591 796 3599 797
rect 2305 769 2357 790
rect 2389 790 3599 796
rect 3651 790 3670 799
rect 3722 790 3741 799
rect 3793 790 3811 799
rect 3863 790 3881 799
rect 3933 790 3951 799
rect 2389 756 2401 790
rect 2435 756 2475 790
rect 2509 756 2549 790
rect 2583 756 2623 790
rect 2657 756 2697 790
rect 2731 756 2771 790
rect 2805 756 2845 790
rect 2879 756 2919 790
rect 2953 756 2993 790
rect 3027 756 3067 790
rect 3101 756 3141 790
rect 3175 756 3215 790
rect 3249 756 3289 790
rect 3323 756 3363 790
rect 3397 756 3437 790
rect 3471 756 3510 790
rect 3544 756 3583 790
rect 3651 756 3656 790
rect 3722 756 3729 790
rect 3793 756 3802 790
rect 3863 756 3875 790
rect 3933 756 3948 790
rect 2389 750 3599 756
tri 3590 747 3593 750 ne
rect 3593 747 3599 750
rect 3651 747 3670 756
rect 3722 747 3741 756
rect 3793 747 3811 756
rect 3863 747 3881 756
rect 3933 747 3951 756
rect 4003 747 4021 799
rect 4073 747 4091 799
rect 4143 747 4161 799
rect 4213 747 4231 799
rect 4283 747 4301 799
rect 4353 747 4359 799
rect 4533 747 4539 799
rect 4591 747 4609 799
rect 4661 747 4679 799
rect 4731 747 4749 799
rect 4801 747 4819 799
rect 4871 747 4889 799
rect 4941 790 4959 799
rect 5011 790 5029 799
rect 5081 790 5099 799
rect 5151 790 5170 799
rect 5222 790 5241 799
rect 5293 790 6162 799
rect 6214 790 6250 799
rect 6302 790 6338 799
rect 6390 790 6503 799
rect 4944 756 4959 790
rect 5017 756 5029 790
rect 5090 756 5099 790
rect 5163 756 5170 790
rect 5236 756 5241 790
rect 5309 756 5348 790
rect 5382 756 5421 790
rect 5455 756 5495 790
rect 5529 756 5569 790
rect 5603 756 5643 790
rect 5677 756 5717 790
rect 5751 756 5791 790
rect 5825 756 5865 790
rect 5899 756 5939 790
rect 5973 756 6013 790
rect 6047 756 6087 790
rect 6121 756 6161 790
rect 6214 756 6235 790
rect 6302 756 6309 790
rect 6417 756 6457 790
rect 6491 756 6503 790
rect 4941 747 4959 756
rect 5011 747 5029 756
rect 5081 747 5099 756
rect 5151 747 5170 756
rect 5222 747 5241 756
rect 5293 747 6162 756
rect 6214 747 6250 756
rect 6302 747 6338 756
rect 6390 747 6503 756
rect 6541 764 6587 803
rect 2305 697 2357 717
rect 6541 730 6547 764
rect 6581 730 6587 764
rect 6541 710 6587 730
rect 6621 1127 6627 1161
rect 6661 1127 6699 1161
rect 6733 1127 6840 1161
rect 6621 1088 6840 1127
rect 6621 1054 6627 1088
rect 6661 1054 6699 1088
rect 6733 1054 6840 1088
rect 6621 1015 6840 1054
rect 6621 981 6627 1015
rect 6661 981 6699 1015
rect 6733 981 6840 1015
rect 6621 942 6840 981
rect 6621 908 6627 942
rect 6661 908 6699 942
rect 6733 908 6840 942
rect 6621 869 6840 908
rect 6621 835 6627 869
rect 6661 835 6699 869
rect 6733 835 6840 869
rect 6621 796 6840 835
rect 6621 762 6627 796
rect 6661 762 6699 796
rect 6733 762 6840 796
rect 6621 723 6840 762
rect 2305 639 2357 645
rect 6539 704 6591 710
tri 3127 640 3130 643 se
rect 3130 640 3136 643
rect 2389 634 3136 640
rect 2153 600 2271 614
tri 2271 600 2304 633 sw
rect 2389 600 2401 634
rect 2435 600 2475 634
rect 2509 600 2549 634
rect 2583 600 2623 634
rect 2657 600 2697 634
rect 2731 600 2771 634
rect 2805 600 2845 634
rect 2879 600 2919 634
rect 2953 600 2993 634
rect 3027 600 3067 634
rect 3101 600 3136 634
rect 2153 594 2304 600
tri 2304 594 2310 600 sw
rect 2389 594 3136 600
rect 2153 579 2310 594
tri 2310 579 2325 594 sw
tri 3127 591 3130 594 ne
rect 3130 591 3136 594
rect 3188 591 3203 643
rect 3255 591 3269 643
rect 3321 634 3335 643
rect 3387 634 3401 643
rect 3453 640 3459 643
tri 3459 640 3462 643 sw
rect 3453 634 4359 640
rect 3323 600 3335 634
rect 3397 600 3401 634
rect 3471 600 3510 634
rect 3544 600 3583 634
rect 3617 600 3656 634
rect 3690 600 3729 634
rect 3763 600 3802 634
rect 3836 600 3875 634
rect 3909 600 3948 634
rect 3982 600 4021 634
rect 4055 600 4094 634
rect 4128 600 4167 634
rect 4201 600 4240 634
rect 4274 600 4313 634
rect 4347 600 4359 634
rect 3321 591 3335 600
rect 3387 591 3401 600
rect 3453 594 4359 600
rect 4533 634 5820 643
rect 5872 634 5885 643
rect 5937 634 5949 643
rect 4533 600 4545 634
rect 4579 600 4618 634
rect 4652 600 4691 634
rect 4725 600 4764 634
rect 4798 600 4837 634
rect 4871 600 4910 634
rect 4944 600 4983 634
rect 5017 600 5056 634
rect 5090 600 5129 634
rect 5163 600 5202 634
rect 5236 600 5275 634
rect 5309 600 5348 634
rect 5382 600 5421 634
rect 5455 600 5495 634
rect 5529 600 5569 634
rect 5603 600 5643 634
rect 5677 600 5717 634
rect 5751 600 5791 634
rect 5937 600 5939 634
rect 3453 591 3459 594
tri 3459 591 3462 594 nw
rect 4533 591 5820 600
rect 5872 591 5885 600
rect 5937 591 5949 600
rect 6001 591 6013 643
rect 6065 591 6077 643
rect 6129 591 6141 643
rect 6193 634 6205 643
rect 6257 634 6269 643
rect 6321 634 6333 643
rect 6385 634 6397 643
rect 6449 634 6503 643
rect 6195 600 6205 634
rect 6449 600 6457 634
rect 6491 600 6503 634
rect 6193 591 6205 600
rect 6257 591 6269 600
rect 6321 591 6333 600
rect 6385 591 6397 600
rect 6449 591 6503 600
rect 6539 631 6591 652
rect 2153 577 2325 579
tri 2325 577 2327 579 sw
rect 2153 575 2327 577
rect 2153 541 2159 575
rect 2193 541 2231 575
rect 2265 573 2327 575
tri 2327 573 2331 577 sw
rect 6539 573 6591 579
rect 6621 689 6627 723
rect 6661 689 6699 723
rect 6733 689 6840 723
rect 6621 650 6840 689
rect 6621 616 6627 650
rect 6661 616 6699 650
rect 6733 616 6840 650
rect 6621 577 6840 616
rect 2265 559 2331 573
tri 2331 559 2345 573 sw
rect 2265 543 2345 559
tri 2345 543 2361 559 sw
tri 6605 543 6621 559 se
rect 6621 543 6627 577
rect 6661 543 6699 577
rect 6733 543 6840 577
rect 2265 541 2361 543
tri 2361 541 2363 543 sw
tri 6603 541 6605 543 se
rect 6605 541 6840 543
rect 2153 539 2363 541
tri 2363 539 2365 541 sw
tri 6601 539 6603 541 se
rect 6603 539 6840 541
rect 2153 505 2365 539
tri 2365 505 2399 539 sw
tri 6567 505 6601 539 se
rect 6601 505 6840 539
rect 2153 504 2399 505
tri 2399 504 2400 505 sw
tri 6566 504 6567 505 se
rect 6567 504 6840 505
rect 2153 502 2400 504
rect 2153 324 2159 502
rect 2265 487 2400 502
tri 2400 487 2417 504 sw
tri 6549 487 6566 504 se
rect 6566 487 6627 504
rect 2265 478 3599 487
rect 3651 478 3670 487
rect 3722 478 3741 487
rect 3793 478 3811 487
rect 3863 478 3881 487
rect 3933 478 3951 487
rect 2265 444 2401 478
rect 2435 444 2475 478
rect 2509 444 2549 478
rect 2583 444 2623 478
rect 2657 444 2697 478
rect 2731 444 2771 478
rect 2805 444 2845 478
rect 2879 444 2919 478
rect 2953 444 2993 478
rect 3027 444 3067 478
rect 3101 444 3141 478
rect 3175 444 3215 478
rect 3249 444 3289 478
rect 3323 444 3363 478
rect 3397 444 3437 478
rect 3471 444 3510 478
rect 3544 444 3583 478
rect 3651 444 3656 478
rect 3722 444 3729 478
rect 3793 444 3802 478
rect 3863 444 3875 478
rect 3933 444 3948 478
rect 2265 435 3599 444
rect 3651 435 3670 444
rect 3722 435 3741 444
rect 3793 435 3811 444
rect 3863 435 3881 444
rect 3933 435 3951 444
rect 4003 435 4021 487
rect 4073 435 4091 487
rect 4143 435 4161 487
rect 4213 435 4231 487
rect 4283 435 4301 487
rect 4353 435 4539 487
rect 4591 435 4609 487
rect 4661 435 4679 487
rect 4731 435 4749 487
rect 4801 435 4819 487
rect 4871 435 4889 487
rect 4941 478 4959 487
rect 5011 478 5029 487
rect 5081 478 5099 487
rect 5151 478 5170 487
rect 5222 478 5241 487
rect 5293 478 6627 487
rect 4944 444 4959 478
rect 5017 444 5029 478
rect 5090 444 5099 478
rect 5163 444 5170 478
rect 5236 444 5241 478
rect 5309 444 5348 478
rect 5382 444 5421 478
rect 5455 444 5495 478
rect 5529 444 5569 478
rect 5603 444 5643 478
rect 5677 444 5717 478
rect 5751 444 5791 478
rect 5825 444 5865 478
rect 5899 444 5939 478
rect 5973 444 6013 478
rect 6047 444 6087 478
rect 6121 444 6161 478
rect 6195 456 6235 478
rect 6269 456 6309 478
rect 6343 456 6383 478
rect 6363 444 6383 456
rect 6417 444 6457 478
rect 6491 470 6627 478
rect 6661 470 6699 504
rect 6733 470 6840 504
rect 6491 444 6840 470
rect 4941 435 4959 444
rect 5011 435 5029 444
rect 5081 435 5099 444
rect 5151 435 5170 444
rect 5222 435 5241 444
rect 5293 435 6183 444
rect 2265 414 6183 435
rect 2265 362 3599 414
rect 3651 362 3665 414
rect 3717 362 3731 414
rect 3783 362 3797 414
rect 3849 362 3863 414
rect 3915 362 3929 414
rect 3981 362 3995 414
rect 4047 362 4061 414
rect 4113 362 4127 414
rect 4179 362 4193 414
rect 4245 362 4259 414
rect 4311 362 4325 414
rect 4377 362 4391 414
rect 4443 362 4457 414
rect 4509 362 4523 414
rect 4575 362 4589 414
rect 4641 362 4655 414
rect 4707 362 4721 414
rect 4773 362 4786 414
rect 4838 362 4851 414
rect 4903 362 4916 414
rect 4968 362 4981 414
rect 5033 362 5046 414
rect 5098 362 5111 414
rect 5163 362 5176 414
rect 5228 362 5241 414
rect 5293 362 6183 414
rect 2265 358 6183 362
rect 6363 431 6840 444
rect 6363 397 6627 431
rect 6661 397 6699 431
rect 6733 397 6840 431
rect 6363 358 6840 397
rect 2265 324 2304 358
rect 2338 324 2377 358
rect 2411 324 2450 358
rect 2484 324 2523 358
rect 2153 286 2523 324
rect 2153 252 2231 286
rect 2265 252 2304 286
rect 2338 252 2377 286
rect 2411 252 2450 286
rect 2484 252 2523 286
rect 6661 324 6699 358
rect 6733 324 6840 358
rect 6661 252 6840 324
rect 2153 246 6840 252
rect 6876 1416 6994 1618
rect 6876 1382 6882 1416
rect 6916 1382 6954 1416
rect 6988 1382 6994 1416
rect 6876 1343 6994 1382
rect 6876 1309 6882 1343
rect 6916 1309 6954 1343
rect 6988 1309 6994 1343
rect 6876 1270 6994 1309
rect 6876 1236 6882 1270
rect 6916 1236 6954 1270
rect 6988 1236 6994 1270
rect 6876 1197 6994 1236
rect 6876 1163 6882 1197
rect 6916 1163 6954 1197
rect 6988 1163 6994 1197
rect 6876 1124 6994 1163
rect 6876 1090 6882 1124
rect 6916 1090 6954 1124
rect 6988 1090 6994 1124
rect 6876 1051 6994 1090
rect 6876 1017 6882 1051
rect 6916 1017 6954 1051
rect 6988 1017 6994 1051
rect 6876 978 6994 1017
rect 6876 944 6882 978
rect 6916 944 6954 978
rect 6988 944 6994 978
rect 6876 905 6994 944
rect 6876 871 6882 905
rect 6916 871 6954 905
rect 6988 871 6994 905
rect 6876 832 6994 871
rect 6876 798 6882 832
rect 6916 798 6954 832
rect 6988 798 6994 832
rect 6876 759 6994 798
rect 6876 725 6882 759
rect 6916 725 6954 759
rect 6988 725 6994 759
rect 6876 686 6994 725
rect 6876 652 6882 686
rect 6916 652 6954 686
rect 6988 652 6994 686
rect 6876 613 6994 652
rect 6876 579 6882 613
rect 6916 579 6954 613
rect 6988 579 6994 613
rect 6876 539 6994 579
rect 6876 505 6882 539
rect 6916 505 6954 539
rect 6988 505 6994 539
rect 6876 465 6994 505
rect 6876 431 6882 465
rect 6916 431 6954 465
rect 6988 431 6994 465
rect 6876 391 6994 431
rect 6876 357 6882 391
rect 6916 357 6954 391
rect 6988 357 6994 391
rect 6876 317 6994 357
rect 6876 283 6882 317
rect 6916 283 6954 317
rect 6988 283 6994 317
tri 173 209 194 230 sw
tri 1877 209 1898 230 se
rect 1898 209 1904 243
rect 1938 209 1976 243
rect 2010 209 2016 243
rect 6876 243 6994 283
rect 167 177 194 209
tri 194 177 226 209 sw
tri 1845 177 1877 209 se
rect 1877 177 2016 209
tri 2016 177 2069 230 sw
tri 6823 177 6876 230 se
rect 6876 177 6882 243
rect 167 171 6882 177
rect 6988 211 6994 243
rect 7157 1450 8618 1456
rect 8670 1450 8684 1456
rect 8736 1450 8750 1456
rect 8802 1450 8816 1456
rect 8868 1450 8882 1456
rect 8934 1450 8948 1456
rect 9000 1450 9014 1456
rect 9066 1450 9080 1456
rect 9132 1450 9146 1456
rect 9198 1450 9212 1456
rect 9264 1450 9278 1456
rect 9330 1450 9344 1456
rect 9396 1450 9410 1456
rect 9462 1450 9476 1456
rect 9528 1450 9542 1456
rect 9594 1450 9608 1456
rect 9660 1450 9674 1456
rect 9726 1450 9740 1456
rect 9792 1450 9805 1456
rect 9857 1450 9870 1456
rect 9922 1450 9935 1456
rect 9987 1450 10000 1456
rect 10052 1450 10065 1456
rect 10117 1450 10130 1456
rect 10182 1450 10195 1456
rect 10247 1450 10260 1456
rect 10312 1450 11757 1456
rect 7157 1416 7241 1450
rect 7275 1416 7319 1450
rect 7353 1416 7397 1450
rect 7431 1416 7475 1450
rect 7509 1416 7553 1450
rect 7587 1416 7631 1450
rect 7665 1416 7709 1450
rect 7743 1416 7788 1450
rect 7822 1416 7898 1450
rect 7157 1378 7898 1416
rect 11460 1416 11499 1450
rect 11533 1416 11572 1450
rect 11606 1416 11645 1450
rect 11679 1416 11757 1450
rect 7157 1344 7163 1378
rect 7197 1344 7235 1378
rect 7269 1344 7319 1378
rect 7353 1344 7397 1378
rect 7431 1344 7475 1378
rect 7509 1344 7553 1378
rect 7587 1344 7631 1378
rect 7665 1344 7709 1378
rect 7743 1344 7788 1378
rect 7822 1344 7898 1378
rect 11460 1378 11757 1416
rect 11460 1344 11499 1378
rect 11533 1344 11572 1378
rect 11606 1344 11645 1378
rect 7157 1340 8618 1344
rect 8670 1340 8684 1344
rect 8736 1340 8750 1344
rect 8802 1340 8816 1344
rect 8868 1340 8882 1344
rect 8934 1340 8948 1344
rect 9000 1340 9014 1344
rect 9066 1340 9080 1344
rect 9132 1340 9146 1344
rect 9198 1340 9212 1344
rect 9264 1340 9278 1344
rect 9330 1340 9344 1344
rect 9396 1340 9410 1344
rect 9462 1340 9476 1344
rect 9528 1340 9542 1344
rect 9594 1340 9608 1344
rect 9660 1340 9674 1344
rect 9726 1340 9740 1344
rect 9792 1340 9805 1344
rect 9857 1340 9870 1344
rect 9922 1340 9935 1344
rect 9987 1340 10000 1344
rect 10052 1340 10065 1344
rect 10117 1340 10130 1344
rect 10182 1340 10195 1344
rect 10247 1340 10260 1344
rect 10312 1340 11645 1344
rect 7157 1338 11645 1340
rect 7157 1305 7275 1338
rect 7157 1271 7163 1305
rect 7197 1271 7235 1305
rect 7269 1271 7275 1305
tri 7275 1298 7315 1338 nw
tri 11599 1298 11639 1338 ne
rect 7157 1232 7275 1271
tri 7415 1264 7418 1267 se
rect 7418 1264 7424 1267
rect 7157 1198 7163 1232
rect 7197 1198 7235 1232
rect 7269 1198 7275 1232
rect 7408 1258 7424 1264
rect 7476 1258 7496 1267
rect 7408 1224 7420 1258
rect 7476 1224 7494 1258
rect 7408 1218 7424 1224
tri 7415 1215 7418 1218 ne
rect 7418 1215 7424 1218
rect 7476 1215 7496 1224
rect 7548 1215 7568 1267
rect 7620 1215 7639 1267
rect 7691 1215 7710 1267
rect 7762 1215 7781 1267
rect 7833 1215 7852 1267
rect 7904 1215 7923 1267
rect 7975 1215 7994 1267
rect 8046 1264 8059 1267
tri 8059 1264 8062 1267 sw
tri 10449 1264 10452 1267 se
rect 10452 1264 10458 1267
rect 8046 1258 9378 1264
rect 8046 1224 8086 1258
rect 8120 1224 8160 1258
rect 8194 1224 8234 1258
rect 8268 1224 8308 1258
rect 8342 1224 8382 1258
rect 8416 1224 8456 1258
rect 8490 1224 8529 1258
rect 8563 1224 8602 1258
rect 8636 1224 8675 1258
rect 8709 1224 8748 1258
rect 8782 1224 8821 1258
rect 8855 1224 8894 1258
rect 8928 1224 8967 1258
rect 9001 1224 9040 1258
rect 9074 1224 9113 1258
rect 9147 1224 9186 1258
rect 9220 1224 9259 1258
rect 9293 1224 9332 1258
rect 9366 1224 9378 1258
rect 8046 1218 9378 1224
rect 9552 1258 10458 1264
rect 10510 1258 10525 1267
rect 10577 1258 10591 1267
rect 9552 1224 9564 1258
rect 9598 1224 9637 1258
rect 9671 1224 9710 1258
rect 9744 1224 9783 1258
rect 9817 1224 9856 1258
rect 9890 1224 9929 1258
rect 9963 1224 10002 1258
rect 10036 1224 10075 1258
rect 10109 1224 10148 1258
rect 10182 1224 10221 1258
rect 10255 1224 10294 1258
rect 10328 1224 10367 1258
rect 10401 1224 10440 1258
rect 10510 1224 10514 1258
rect 10577 1224 10588 1258
rect 9552 1218 10458 1224
rect 8046 1215 8059 1218
tri 8059 1215 8062 1218 nw
tri 10449 1215 10452 1218 ne
rect 10452 1215 10458 1218
rect 10510 1215 10525 1224
rect 10577 1215 10591 1224
rect 10643 1215 10657 1267
rect 10709 1215 10723 1267
rect 10775 1264 10781 1267
tri 10781 1264 10784 1267 sw
rect 10775 1258 11522 1264
rect 10775 1224 10810 1258
rect 10844 1224 10884 1258
rect 10918 1224 10958 1258
rect 10992 1224 11032 1258
rect 11066 1224 11106 1258
rect 11140 1224 11180 1258
rect 11214 1224 11254 1258
rect 11288 1224 11328 1258
rect 11362 1224 11402 1258
rect 11436 1224 11476 1258
rect 11510 1224 11522 1258
rect 10775 1218 11522 1224
rect 10775 1215 10781 1218
tri 10781 1215 10784 1218 nw
rect 7157 1159 7275 1198
rect 7157 1125 7163 1159
rect 7197 1125 7235 1159
rect 7269 1125 7275 1159
rect 7157 1086 7275 1125
rect 7157 1052 7163 1086
rect 7197 1052 7235 1086
rect 7269 1052 7275 1086
rect 7157 1013 7275 1052
rect 7157 979 7163 1013
rect 7197 979 7235 1013
rect 7269 979 7275 1013
rect 7157 940 7275 979
rect 7157 906 7163 940
rect 7197 906 7235 940
rect 7269 906 7275 940
rect 7157 867 7275 906
rect 7157 833 7163 867
rect 7197 833 7235 867
rect 7269 833 7275 867
rect 7157 794 7275 833
rect 7157 760 7163 794
rect 7197 760 7235 794
rect 7269 760 7275 794
rect 7157 721 7275 760
rect 7157 687 7163 721
rect 7197 687 7235 721
rect 7269 687 7275 721
rect 7157 648 7275 687
rect 7157 614 7163 648
rect 7197 614 7235 648
rect 7269 614 7275 648
rect 7157 575 7275 614
rect 7157 541 7163 575
rect 7197 541 7235 575
rect 7269 541 7275 575
rect 7157 502 7275 541
rect 7157 272 7163 502
rect 7269 397 7275 502
rect 7322 1207 7374 1213
rect 7322 1141 7374 1155
rect 11558 1207 11610 1213
rect 11558 1141 11610 1155
tri 8609 1108 8612 1111 se
rect 8612 1108 8618 1111
rect 7322 1075 7374 1089
rect 7408 1102 8618 1108
rect 8670 1102 8689 1111
rect 8741 1102 8760 1111
rect 8812 1102 8830 1111
rect 8882 1102 8900 1111
rect 8952 1102 8970 1111
rect 7408 1068 7420 1102
rect 7454 1068 7494 1102
rect 7528 1068 7568 1102
rect 7602 1068 7642 1102
rect 7676 1068 7716 1102
rect 7750 1068 7790 1102
rect 7824 1068 7864 1102
rect 7898 1068 7938 1102
rect 7972 1068 8012 1102
rect 8046 1068 8086 1102
rect 8120 1068 8160 1102
rect 8194 1068 8234 1102
rect 8268 1068 8308 1102
rect 8342 1068 8382 1102
rect 8416 1068 8456 1102
rect 8490 1068 8529 1102
rect 8563 1068 8602 1102
rect 8670 1068 8675 1102
rect 8741 1068 8748 1102
rect 8812 1068 8821 1102
rect 8882 1068 8894 1102
rect 8952 1068 8967 1102
rect 7408 1062 8618 1068
tri 8609 1059 8612 1062 ne
rect 8612 1059 8618 1062
rect 8670 1059 8689 1068
rect 8741 1059 8760 1068
rect 8812 1059 8830 1068
rect 8882 1059 8900 1068
rect 8952 1059 8970 1068
rect 9022 1059 9040 1111
rect 9092 1059 9110 1111
rect 9162 1059 9180 1111
rect 9232 1059 9250 1111
rect 9302 1059 9320 1111
rect 9372 1059 9378 1111
rect 9552 1059 9558 1111
rect 9610 1059 9628 1111
rect 9680 1059 9698 1111
rect 9750 1059 9768 1111
rect 9820 1059 9838 1111
rect 9890 1059 9908 1111
rect 9960 1102 9978 1111
rect 10030 1102 10048 1111
rect 10100 1102 10118 1111
rect 10170 1102 10189 1111
rect 10241 1102 10260 1111
rect 10312 1108 10318 1111
tri 10318 1108 10321 1111 sw
rect 10312 1102 11522 1108
rect 9963 1068 9978 1102
rect 10036 1068 10048 1102
rect 10109 1068 10118 1102
rect 10182 1068 10189 1102
rect 10255 1068 10260 1102
rect 10328 1068 10367 1102
rect 10401 1068 10440 1102
rect 10474 1068 10514 1102
rect 10548 1068 10588 1102
rect 10622 1068 10662 1102
rect 10696 1068 10736 1102
rect 10770 1068 10810 1102
rect 10844 1068 10884 1102
rect 10918 1068 10958 1102
rect 10992 1068 11032 1102
rect 11066 1068 11106 1102
rect 11140 1068 11180 1102
rect 11214 1068 11254 1102
rect 11288 1068 11328 1102
rect 11362 1068 11402 1102
rect 11436 1068 11476 1102
rect 11510 1068 11522 1102
rect 9960 1059 9978 1068
rect 10030 1059 10048 1068
rect 10100 1059 10118 1068
rect 10170 1059 10189 1068
rect 10241 1059 10260 1068
rect 10312 1062 11522 1068
rect 11558 1075 11610 1089
rect 10312 1059 10318 1062
tri 10318 1059 10321 1062 nw
rect 7322 1019 7330 1023
rect 7364 1019 7374 1023
rect 7322 1009 7374 1019
rect 7322 945 7330 957
rect 7364 945 7374 957
rect 11558 1019 11566 1023
rect 11600 1019 11610 1023
rect 11558 1009 11610 1019
tri 7415 952 7418 955 se
rect 7418 952 7424 955
rect 7322 943 7374 945
rect 7408 946 7424 952
rect 7476 946 7495 955
rect 7408 912 7420 946
rect 7476 912 7494 946
rect 7408 906 7424 912
tri 7415 905 7416 906 ne
rect 7416 905 7424 906
tri 7416 903 7418 905 ne
rect 7418 903 7424 905
rect 7476 903 7495 912
rect 7547 903 7566 955
rect 7618 903 7637 955
rect 7689 903 7707 955
rect 7759 903 7777 955
rect 7829 903 7847 955
rect 7899 903 7917 955
rect 7969 946 7987 955
rect 8039 952 8045 955
tri 8045 952 8048 955 sw
tri 10449 952 10452 955 se
rect 10452 952 10458 955
rect 8039 946 9378 952
rect 7972 912 7987 946
rect 8046 912 8086 946
rect 8120 912 8160 946
rect 8194 912 8234 946
rect 8268 912 8308 946
rect 8342 912 8382 946
rect 8416 912 8456 946
rect 8490 912 8529 946
rect 8563 912 8602 946
rect 8636 912 8675 946
rect 8709 912 8748 946
rect 8782 912 8821 946
rect 8855 912 8894 946
rect 8928 912 8967 946
rect 9001 912 9040 946
rect 9074 912 9113 946
rect 9147 912 9186 946
rect 9220 912 9259 946
rect 9293 912 9332 946
rect 9366 912 9378 946
rect 7969 903 7987 912
rect 8039 906 9378 912
rect 9552 946 10458 952
rect 10510 946 10525 955
rect 10577 946 10591 955
rect 9552 912 9564 946
rect 9598 912 9637 946
rect 9671 912 9710 946
rect 9744 912 9783 946
rect 9817 912 9856 946
rect 9890 912 9929 946
rect 9963 912 10002 946
rect 10036 912 10075 946
rect 10109 912 10148 946
rect 10182 912 10221 946
rect 10255 912 10294 946
rect 10328 912 10367 946
rect 10401 912 10440 946
rect 10510 912 10514 946
rect 10577 912 10588 946
rect 9552 906 10458 912
rect 8039 905 8047 906
tri 8047 905 8048 906 nw
tri 10449 905 10450 906 ne
rect 10450 905 10458 906
rect 8039 903 8045 905
tri 8045 903 8047 905 nw
tri 10450 903 10452 905 ne
rect 10452 903 10458 905
rect 10510 903 10525 912
rect 10577 903 10591 912
rect 10643 903 10657 955
rect 10709 903 10723 955
rect 10775 952 10781 955
tri 10781 952 10784 955 sw
rect 10775 946 11522 952
rect 10775 912 10810 946
rect 10844 912 10884 946
rect 10918 912 10958 946
rect 10992 912 11032 946
rect 11066 912 11106 946
rect 11140 912 11180 946
rect 11214 912 11254 946
rect 11288 912 11328 946
rect 11362 912 11402 946
rect 11436 912 11476 946
rect 11510 912 11522 946
rect 10775 906 11522 912
rect 11558 945 11566 957
rect 11600 945 11610 957
rect 11558 943 11610 945
rect 10775 905 10783 906
tri 10783 905 10784 906 nw
rect 10775 903 10781 905
tri 10781 903 10783 905 nw
rect 7322 877 7330 891
rect 7364 877 7374 891
rect 7322 811 7330 825
rect 7364 811 7374 825
rect 11558 877 11566 891
rect 11600 877 11610 891
rect 11558 811 11566 825
rect 11600 811 11610 825
tri 8610 797 8612 799 se
rect 8612 797 8618 799
tri 8609 796 8610 797 se
rect 8610 796 8618 797
rect 7322 757 7374 759
rect 7322 745 7330 757
rect 7364 745 7374 757
rect 7408 790 8618 796
rect 8670 790 8689 799
rect 8741 790 8760 799
rect 8812 790 8830 799
rect 8882 790 8900 799
rect 8952 790 8970 799
rect 7408 756 7420 790
rect 7454 756 7494 790
rect 7528 756 7568 790
rect 7602 756 7642 790
rect 7676 756 7716 790
rect 7750 756 7790 790
rect 7824 756 7864 790
rect 7898 756 7938 790
rect 7972 756 8012 790
rect 8046 756 8086 790
rect 8120 756 8160 790
rect 8194 756 8234 790
rect 8268 756 8308 790
rect 8342 756 8382 790
rect 8416 756 8456 790
rect 8490 756 8529 790
rect 8563 756 8602 790
rect 8670 756 8675 790
rect 8741 756 8748 790
rect 8812 756 8821 790
rect 8882 756 8894 790
rect 8952 756 8967 790
rect 7408 750 8618 756
tri 8609 747 8612 750 ne
rect 8612 747 8618 750
rect 8670 747 8689 756
rect 8741 747 8760 756
rect 8812 747 8830 756
rect 8882 747 8900 756
rect 8952 747 8970 756
rect 9022 747 9040 799
rect 9092 747 9110 799
rect 9162 747 9180 799
rect 9232 747 9250 799
rect 9302 747 9320 799
rect 9372 747 9378 799
rect 9552 747 9558 799
rect 9610 747 9628 799
rect 9680 747 9698 799
rect 9750 747 9768 799
rect 9820 747 9838 799
rect 9890 747 9908 799
rect 9960 790 9978 799
rect 10030 790 10048 799
rect 10100 790 10118 799
rect 10170 790 10189 799
rect 10241 790 10260 799
rect 10312 797 10318 799
tri 10318 797 10320 799 sw
rect 10312 796 10320 797
tri 10320 796 10321 797 sw
rect 10312 790 11522 796
rect 9963 756 9978 790
rect 10036 756 10048 790
rect 10109 756 10118 790
rect 10182 756 10189 790
rect 10255 756 10260 790
rect 10328 756 10367 790
rect 10401 756 10440 790
rect 10474 756 10514 790
rect 10548 756 10588 790
rect 10622 756 10662 790
rect 10696 756 10736 790
rect 10770 756 10810 790
rect 10844 756 10884 790
rect 10918 756 10958 790
rect 10992 756 11032 790
rect 11066 756 11106 790
rect 11140 756 11180 790
rect 11214 756 11254 790
rect 11288 756 11328 790
rect 11362 756 11402 790
rect 11436 756 11476 790
rect 11510 756 11522 790
rect 9960 747 9978 756
rect 10030 747 10048 756
rect 10100 747 10118 756
rect 10170 747 10189 756
rect 10241 747 10260 756
rect 10312 750 11522 756
rect 11558 757 11610 759
rect 10312 747 10318 750
tri 10318 747 10321 750 nw
rect 7322 683 7374 693
rect 7322 679 7330 683
rect 7364 679 7374 683
rect 11558 745 11566 757
rect 11600 745 11610 757
rect 11558 683 11610 693
rect 11558 679 11566 683
rect 11600 679 11610 683
tri 7415 640 7418 643 se
rect 7418 640 7424 643
rect 7322 613 7374 627
rect 7408 634 7424 640
rect 7476 634 7496 643
rect 7408 600 7420 634
rect 7476 600 7494 634
rect 7408 594 7424 600
tri 7415 591 7418 594 ne
rect 7418 591 7424 594
rect 7476 591 7496 600
rect 7548 591 7568 643
rect 7620 591 7639 643
rect 7691 591 7710 643
rect 7762 591 7781 643
rect 7833 591 7852 643
rect 7904 591 7923 643
rect 7975 591 7994 643
rect 8046 640 8052 643
tri 8052 640 8055 643 sw
tri 10449 640 10452 643 se
rect 10452 640 10458 643
rect 8046 634 9378 640
rect 8046 600 8086 634
rect 8120 600 8160 634
rect 8194 600 8234 634
rect 8268 600 8308 634
rect 8342 600 8382 634
rect 8416 600 8456 634
rect 8490 600 8529 634
rect 8563 600 8602 634
rect 8636 600 8675 634
rect 8709 600 8748 634
rect 8782 600 8821 634
rect 8855 600 8894 634
rect 8928 600 8967 634
rect 9001 600 9040 634
rect 9074 600 9113 634
rect 9147 600 9186 634
rect 9220 600 9259 634
rect 9293 600 9332 634
rect 9366 600 9378 634
rect 8046 594 9378 600
rect 9552 634 10458 640
rect 10510 634 10525 643
rect 10577 634 10591 643
rect 9552 600 9564 634
rect 9598 600 9637 634
rect 9671 600 9710 634
rect 9744 600 9783 634
rect 9817 600 9856 634
rect 9890 600 9929 634
rect 9963 600 10002 634
rect 10036 600 10075 634
rect 10109 600 10148 634
rect 10182 600 10221 634
rect 10255 600 10294 634
rect 10328 600 10367 634
rect 10401 600 10440 634
rect 10510 600 10514 634
rect 10577 600 10588 634
rect 9552 594 10458 600
rect 8046 591 8052 594
tri 8052 591 8055 594 nw
tri 10449 591 10452 594 ne
rect 10452 591 10458 594
rect 10510 591 10525 600
rect 10577 591 10591 600
rect 10643 591 10657 643
rect 10709 591 10723 643
rect 10775 640 10781 643
tri 10781 640 10784 643 sw
rect 10775 634 11522 640
rect 10775 600 10810 634
rect 10844 600 10884 634
rect 10918 600 10958 634
rect 10992 600 11032 634
rect 11066 600 11106 634
rect 11140 600 11180 634
rect 11214 600 11254 634
rect 11288 600 11328 634
rect 11362 600 11402 634
rect 11436 600 11476 634
rect 11510 600 11522 634
rect 10775 594 11522 600
rect 11558 613 11610 627
rect 10775 591 10781 594
tri 10781 591 10784 594 nw
rect 7322 547 7374 561
rect 7322 489 7374 495
rect 11558 547 11610 561
rect 11558 489 11610 495
rect 11639 1200 11645 1338
rect 11751 1200 11757 1378
rect 11639 1161 11757 1200
rect 11639 1127 11645 1161
rect 11679 1127 11717 1161
rect 11751 1127 11757 1161
rect 11639 1088 11757 1127
rect 11639 1054 11645 1088
rect 11679 1054 11717 1088
rect 11751 1054 11757 1088
rect 11639 1015 11757 1054
rect 11639 981 11645 1015
rect 11679 981 11717 1015
rect 11751 981 11757 1015
rect 11639 942 11757 981
rect 11639 908 11645 942
rect 11679 908 11717 942
rect 11751 908 11757 942
rect 11639 869 11757 908
rect 11639 835 11645 869
rect 11679 835 11717 869
rect 11751 835 11757 869
rect 11639 796 11757 835
rect 11639 762 11645 796
rect 11679 762 11717 796
rect 11751 762 11757 796
rect 11639 723 11757 762
rect 11639 689 11645 723
rect 11679 689 11717 723
rect 11751 689 11757 723
rect 11639 650 11757 689
rect 11639 616 11645 650
rect 11679 616 11717 650
rect 11751 616 11757 650
rect 11639 577 11757 616
rect 11639 543 11645 577
rect 11679 543 11717 577
rect 11751 543 11757 577
rect 11639 504 11757 543
tri 8609 484 8612 487 se
rect 8612 484 8618 487
rect 7408 478 8618 484
rect 8670 478 8689 487
rect 8741 478 8760 487
rect 8812 478 8830 487
rect 8882 478 8900 487
rect 8952 478 8970 487
rect 7408 444 7420 478
rect 7454 444 7494 478
rect 7528 444 7568 478
rect 7602 444 7642 478
rect 7676 444 7716 478
rect 7750 444 7790 478
rect 7824 444 7864 478
rect 7898 444 7938 478
rect 7972 444 8012 478
rect 8046 444 8086 478
rect 8120 444 8160 478
rect 8194 444 8234 478
rect 8268 444 8308 478
rect 8342 444 8382 478
rect 8416 444 8456 478
rect 8490 444 8529 478
rect 8563 444 8602 478
rect 8670 444 8675 478
rect 8741 444 8748 478
rect 8812 444 8821 478
rect 8882 444 8894 478
rect 8952 444 8967 478
rect 7408 438 8618 444
tri 8609 435 8612 438 ne
rect 8612 435 8618 438
rect 8670 435 8689 444
rect 8741 435 8760 444
rect 8812 435 8830 444
rect 8882 435 8900 444
rect 8952 435 8970 444
rect 9022 435 9040 487
rect 9092 435 9110 487
rect 9162 435 9180 487
rect 9232 435 9250 487
rect 9302 435 9320 487
rect 9372 435 9378 487
rect 9552 435 9558 487
rect 9610 435 9628 487
rect 9680 435 9698 487
rect 9750 435 9768 487
rect 9820 435 9838 487
rect 9890 435 9908 487
rect 9960 478 9978 487
rect 10030 478 10048 487
rect 10100 478 10118 487
rect 10170 478 10189 487
rect 10241 478 10260 487
rect 10312 484 10318 487
tri 10318 484 10321 487 sw
rect 10312 478 11522 484
rect 9963 444 9978 478
rect 10036 444 10048 478
rect 10109 444 10118 478
rect 10182 444 10189 478
rect 10255 444 10260 478
rect 10328 444 10367 478
rect 10401 444 10440 478
rect 10474 444 10514 478
rect 10548 444 10588 478
rect 10622 444 10662 478
rect 10696 444 10736 478
rect 10770 444 10810 478
rect 10844 444 10884 478
rect 10918 444 10958 478
rect 10992 444 11032 478
rect 11066 444 11106 478
rect 11140 444 11180 478
rect 11214 444 11254 478
rect 11288 444 11328 478
rect 11362 444 11402 478
rect 11436 444 11476 478
rect 11510 444 11522 478
rect 9960 435 9978 444
rect 10030 435 10048 444
rect 10100 435 10118 444
rect 10170 435 10189 444
rect 10241 435 10260 444
rect 10312 438 11522 444
rect 11639 470 11645 504
rect 11679 470 11717 504
rect 11751 470 11757 504
rect 10312 435 10318 438
tri 10318 435 10321 438 nw
rect 11639 431 11757 470
tri 7275 397 7295 417 sw
tri 11619 397 11639 417 se
rect 11639 397 11645 431
rect 11679 397 11717 431
rect 11751 397 11757 431
rect 7269 393 7295 397
tri 7295 393 7299 397 sw
tri 11615 393 11619 397 se
rect 11619 393 11757 397
rect 7269 364 7299 393
tri 7299 364 7328 393 sw
tri 11605 383 11615 393 se
rect 11615 383 11757 393
tri 8593 364 8612 383 se
rect 8612 364 8618 383
rect 7269 358 8618 364
rect 8670 358 8684 383
rect 8736 358 8750 383
rect 8802 358 8816 383
rect 8868 358 8882 383
rect 8934 358 8948 383
rect 9000 358 9014 383
rect 9066 358 9080 383
rect 9132 358 9146 383
rect 9198 358 9212 383
rect 9264 358 9278 383
rect 9330 358 9344 383
rect 9396 358 9410 383
rect 9462 358 9476 383
rect 9528 358 9542 383
rect 9594 358 9608 383
rect 9660 358 9674 383
rect 9726 358 9740 383
rect 9792 358 9805 383
rect 9857 358 9870 383
rect 9922 358 9935 383
rect 9987 358 10000 383
rect 10052 358 10065 383
rect 10117 358 10130 383
rect 10182 358 10195 383
rect 10247 358 10260 383
rect 10312 364 10318 383
tri 10318 364 10337 383 sw
tri 11586 364 11605 383 se
rect 11605 364 11757 383
rect 10312 358 11757 364
rect 7269 324 7308 358
rect 7342 324 7381 358
rect 7415 324 7454 358
rect 7488 324 7527 358
rect 7561 324 7600 358
rect 7634 324 7673 358
rect 7707 324 7746 358
rect 7780 324 7819 358
rect 7853 324 7892 358
rect 7926 324 7965 358
rect 7999 324 8038 358
rect 8072 324 8111 358
rect 8145 324 8184 358
rect 8218 324 8257 358
rect 8291 324 8330 358
rect 8364 324 8403 358
rect 8437 324 8476 358
rect 8510 324 8549 358
rect 7215 272 7229 324
rect 7281 272 7295 324
rect 7347 272 7361 324
rect 7413 286 7426 324
rect 7478 286 7491 324
rect 7543 286 7556 324
rect 7608 286 7621 324
rect 7673 286 7686 324
rect 7738 286 7751 324
rect 7415 272 7426 286
rect 7488 272 7491 286
rect 7738 272 7746 286
rect 7803 272 7816 324
rect 7868 272 7881 324
rect 7933 272 7946 324
rect 7998 286 8011 324
rect 8063 286 8076 324
rect 8128 286 8549 324
rect 11679 324 11717 358
rect 11751 324 11757 358
rect 7999 272 8011 286
rect 8072 272 8076 286
rect 7157 260 7235 272
rect 7269 260 7308 272
rect 7342 260 7381 272
rect 7415 260 7454 272
rect 7488 260 7527 272
rect 7561 260 7600 272
rect 7634 260 7673 272
rect 7707 260 7746 272
rect 7780 260 7819 272
rect 7853 260 7892 272
rect 7926 260 7965 272
rect 7999 260 8038 272
rect 8072 260 8111 272
tri 6994 211 7013 230 sw
rect 6988 208 7013 211
tri 7013 208 7016 211 sw
rect 7157 208 7163 260
rect 7215 208 7229 260
rect 7281 208 7295 260
rect 7347 208 7361 260
rect 7415 252 7426 260
rect 7488 252 7491 260
rect 7738 252 7746 260
rect 7413 208 7426 252
rect 7478 208 7491 252
rect 7543 208 7556 252
rect 7608 208 7621 252
rect 7673 208 7686 252
rect 7738 208 7751 252
rect 7803 208 7816 260
rect 7868 208 7881 260
rect 7933 208 7946 260
rect 7999 252 8011 260
rect 8072 252 8076 260
rect 8145 252 8184 286
rect 8218 252 8257 286
rect 8291 252 8330 286
rect 8364 252 8403 286
rect 8437 252 8476 286
rect 8510 252 8549 286
rect 11679 252 11757 324
rect 7998 208 8011 252
rect 8063 208 8076 252
rect 8128 246 11757 252
rect 11894 1425 12012 1463
rect 11894 1391 11900 1425
rect 11934 1391 11972 1425
rect 12006 1391 12012 1425
rect 11894 1352 12012 1391
rect 11894 1318 11900 1352
rect 11934 1318 11972 1352
rect 12006 1318 12012 1352
rect 11894 1279 12012 1318
rect 11894 1245 11900 1279
rect 11934 1245 11972 1279
rect 12006 1245 12012 1279
rect 11894 1206 12012 1245
rect 11894 1172 11900 1206
rect 11934 1172 11972 1206
rect 12006 1172 12012 1206
rect 11894 1133 12012 1172
rect 11894 1099 11900 1133
rect 11934 1099 11972 1133
rect 12006 1099 12012 1133
rect 11894 1059 12012 1099
rect 11894 1025 11900 1059
rect 11934 1025 11972 1059
rect 12006 1025 12012 1059
rect 11894 985 12012 1025
rect 11894 951 11900 985
rect 11934 951 11972 985
rect 12006 951 12012 985
rect 11894 911 12012 951
rect 11894 877 11900 911
rect 11934 877 11972 911
rect 12006 877 12012 911
rect 11894 837 12012 877
rect 11894 803 11900 837
rect 11934 803 11972 837
rect 12006 803 12012 837
rect 11894 763 12012 803
rect 11894 729 11900 763
rect 11934 729 11972 763
rect 12006 729 12012 763
rect 11894 689 12012 729
rect 11894 655 11900 689
rect 11934 655 11972 689
rect 12006 655 12012 689
rect 11894 615 12012 655
rect 11894 581 11900 615
rect 11934 581 11972 615
rect 12006 581 12012 615
rect 11894 541 12012 581
rect 11894 507 11900 541
rect 11934 507 11972 541
rect 12006 507 12012 541
rect 11894 467 12012 507
rect 11894 433 11900 467
rect 11934 433 11972 467
rect 12006 433 12012 467
rect 11894 393 12012 433
rect 11894 359 11900 393
rect 11934 359 11972 393
rect 12006 359 12012 393
rect 11894 319 12012 359
rect 11894 285 11900 319
rect 11934 285 11972 319
rect 12006 285 12012 319
rect 8128 245 8171 246
tri 8171 245 8172 246 nw
rect 11894 245 12012 285
rect 8128 211 8137 245
tri 8137 211 8171 245 nw
tri 11875 211 11894 230 se
rect 11894 211 11900 245
rect 11934 211 11972 245
rect 12006 211 12012 245
rect 8128 208 8134 211
tri 8134 208 8137 211 nw
tri 11872 208 11875 211 se
rect 11875 208 12012 211
rect 6988 177 7016 208
tri 7016 177 7047 208 sw
tri 11841 177 11872 208 se
rect 11872 177 12012 208
rect 6988 171 12012 177
rect 167 137 206 171
rect 240 137 279 171
rect 313 137 352 171
rect 386 137 425 171
rect 459 137 498 171
rect 532 137 571 171
rect 605 137 644 171
rect 678 137 717 171
rect 751 137 790 171
rect 824 137 863 171
rect 897 137 936 171
rect 970 137 1009 171
rect 1043 137 1082 171
rect 1116 137 1155 171
rect 1189 137 1228 171
rect 1262 137 1301 171
rect 1335 137 1374 171
rect 1408 137 1447 171
rect 1481 137 1520 171
rect 1554 137 1593 171
rect 1627 137 1666 171
rect 1700 137 1739 171
rect 1773 137 1812 171
rect 1846 137 1885 171
rect 1919 137 1958 171
rect 1992 137 2031 171
rect 2065 137 2104 171
rect 2138 137 2177 171
rect 2211 137 2250 171
rect 2284 137 2323 171
rect 2357 137 2396 171
rect 55 99 2396 137
rect 55 65 133 99
rect 167 65 206 99
rect 240 65 279 99
rect 313 65 352 99
rect 386 65 425 99
rect 459 65 498 99
rect 532 65 571 99
rect 605 65 644 99
rect 678 65 717 99
rect 751 65 790 99
rect 824 65 863 99
rect 897 65 936 99
rect 970 65 1009 99
rect 1043 65 1082 99
rect 1116 65 1155 99
rect 1189 65 1228 99
rect 1262 65 1301 99
rect 1335 65 1374 99
rect 1408 65 1447 99
rect 1481 65 1520 99
rect 1554 65 1593 99
rect 1627 65 1666 99
rect 1700 65 1739 99
rect 1773 65 1812 99
rect 1846 65 1885 99
rect 1919 65 1958 99
rect 1992 65 2031 99
rect 2065 65 2104 99
rect 2138 65 2177 99
rect 2211 65 2250 99
rect 2284 65 2323 99
rect 2357 65 2396 99
rect 11934 137 11972 171
rect 12006 137 12012 171
rect 11934 65 12012 137
rect 55 59 12012 65
rect -508 -54 37 -48
rect -508 -88 -496 -54
rect -462 -88 -409 -54
rect -375 -88 -322 -54
rect -288 -88 -236 -54
rect -202 -56 -150 -54
rect -116 -56 37 -54
rect -202 -88 -195 -56
rect -508 -108 -195 -88
rect -143 -108 -131 -88
rect -79 -108 37 -56
rect -508 -124 37 -108
rect -508 -164 -195 -124
rect -143 -164 -131 -124
rect -508 -198 -496 -164
rect -462 -198 -409 -164
rect -375 -198 -322 -164
rect -288 -198 -236 -164
rect -202 -176 -195 -164
rect -79 -176 37 -124
rect -202 -198 -150 -176
rect -116 -198 37 -176
rect -508 -204 37 -198
rect 5371 -281 5377 -229
rect 5429 -281 5441 -229
rect 5493 -281 5499 -229
rect 5411 -1301 5463 -281
rect 5411 -1365 5463 -1353
rect 5411 -1423 5463 -1417
rect 5611 -1153 7982 -1147
rect 5611 -1187 5691 -1153
rect 5725 -1187 5765 -1153
rect 5799 -1187 5839 -1153
rect 5873 -1187 5913 -1153
rect 5947 -1187 5987 -1153
rect 6021 -1187 6062 -1153
rect 6096 -1187 6137 -1153
rect 6171 -1187 6212 -1153
rect 6246 -1187 6287 -1153
rect 6321 -1187 6397 -1153
rect 6431 -1187 6470 -1153
rect 6504 -1187 6543 -1153
rect 6577 -1187 6616 -1153
rect 6650 -1187 6689 -1153
rect 6723 -1187 6762 -1153
rect 6796 -1187 6835 -1153
rect 6869 -1187 6908 -1153
rect 6942 -1187 6982 -1153
rect 7016 -1187 7056 -1153
rect 7090 -1187 7130 -1153
rect 7164 -1187 7204 -1153
rect 7238 -1187 7278 -1153
rect 7312 -1187 7352 -1153
rect 7386 -1187 7426 -1153
rect 7460 -1187 7500 -1153
rect 7534 -1187 7574 -1153
rect 7608 -1187 7648 -1153
rect 7682 -1187 7722 -1153
rect 7756 -1187 7796 -1153
rect 7830 -1187 7870 -1153
rect 7904 -1187 7982 -1153
rect 5611 -1193 7982 -1187
rect 5611 -1225 5657 -1193
rect 5611 -1259 5617 -1225
rect 5651 -1259 5657 -1225
rect 5611 -1304 5657 -1259
rect 7936 -1231 7982 -1193
rect 5611 -1338 5617 -1304
rect 5651 -1338 5657 -1304
rect 5611 -1383 5657 -1338
rect 5611 -1417 5617 -1383
rect 5651 -1417 5657 -1383
rect 5611 -1462 5657 -1417
rect 5723 -1301 5775 -1295
rect 5840 -1313 5846 -1261
rect 5898 -1313 5911 -1261
rect 5963 -1313 5976 -1261
rect 6028 -1270 6041 -1261
rect 6093 -1270 6106 -1261
rect 6158 -1270 6171 -1261
rect 6223 -1270 6236 -1261
rect 6036 -1304 6041 -1270
rect 6223 -1304 6227 -1270
rect 6028 -1313 6041 -1304
rect 6093 -1313 6106 -1304
rect 6158 -1313 6171 -1304
rect 6223 -1313 6236 -1304
rect 6288 -1313 6301 -1261
rect 6353 -1313 6365 -1261
rect 6417 -1313 6429 -1261
rect 6481 -1270 6493 -1261
rect 6545 -1270 6557 -1261
rect 6609 -1270 6621 -1261
rect 6673 -1270 6685 -1261
rect 6486 -1304 6493 -1270
rect 6673 -1304 6676 -1270
rect 6481 -1313 6493 -1304
rect 6545 -1313 6557 -1304
rect 6609 -1313 6621 -1304
rect 6673 -1313 6685 -1304
rect 6737 -1313 6749 -1261
rect 6801 -1313 6813 -1261
rect 6865 -1313 6877 -1261
rect 6929 -1270 6941 -1261
rect 6993 -1270 7005 -1261
rect 7057 -1270 7069 -1261
rect 7121 -1270 7133 -1261
rect 7185 -1270 7197 -1261
rect 6932 -1304 6941 -1270
rect 7185 -1304 7194 -1270
rect 6929 -1313 6941 -1304
rect 6993 -1313 7005 -1304
rect 7057 -1313 7069 -1304
rect 7121 -1313 7133 -1304
rect 7185 -1313 7197 -1304
rect 7249 -1313 7261 -1261
rect 7313 -1313 7325 -1261
rect 7377 -1313 7389 -1261
rect 7441 -1270 7453 -1261
rect 7505 -1270 7517 -1261
rect 7569 -1270 7581 -1261
rect 7633 -1270 7645 -1261
rect 7450 -1304 7453 -1270
rect 7633 -1304 7638 -1270
rect 7441 -1313 7453 -1304
rect 7505 -1313 7517 -1304
rect 7569 -1313 7581 -1304
rect 7633 -1313 7645 -1304
rect 7697 -1313 7709 -1261
rect 7761 -1313 7773 -1261
rect 7825 -1264 7831 -1261
rect 7825 -1310 7832 -1264
rect 7936 -1265 7942 -1231
rect 7976 -1265 7982 -1231
rect 7936 -1309 7982 -1265
rect 7825 -1313 7831 -1310
rect 5723 -1361 5734 -1353
rect 5768 -1361 5775 -1353
rect 5723 -1365 5775 -1361
rect 7936 -1343 7942 -1309
rect 7976 -1343 7982 -1309
rect 7936 -1387 7982 -1343
rect 5723 -1423 5734 -1417
rect 5611 -1496 5617 -1462
rect 5651 -1496 5657 -1462
rect 5611 -1541 5657 -1496
rect 5611 -1575 5617 -1541
rect 5651 -1575 5657 -1541
rect 5611 -1620 5657 -1575
rect 5611 -1654 5617 -1620
rect 5651 -1654 5657 -1620
rect 5611 -1698 5657 -1654
rect 5611 -1732 5617 -1698
rect 5651 -1732 5657 -1698
rect 5611 -1776 5657 -1732
rect 5611 -1810 5617 -1776
rect 5651 -1810 5657 -1776
rect 5611 -1854 5657 -1810
rect 5611 -1888 5617 -1854
rect 5651 -1888 5657 -1854
rect 5728 -1433 5734 -1423
rect 5768 -1423 5775 -1417
rect 5768 -1433 5774 -1423
rect 5728 -1472 5774 -1433
rect 5840 -1469 5846 -1417
rect 5898 -1469 5911 -1417
rect 5963 -1469 5976 -1417
rect 6028 -1426 6041 -1417
rect 6093 -1426 6106 -1417
rect 6158 -1426 6171 -1417
rect 6223 -1426 6236 -1417
rect 6036 -1460 6041 -1426
rect 6223 -1460 6227 -1426
rect 6028 -1469 6041 -1460
rect 6093 -1469 6106 -1460
rect 6158 -1469 6171 -1460
rect 6223 -1469 6236 -1460
rect 6288 -1469 6301 -1417
rect 6353 -1469 6365 -1417
rect 6417 -1469 6429 -1417
rect 6481 -1426 6493 -1417
rect 6545 -1426 6557 -1417
rect 6609 -1426 6621 -1417
rect 6673 -1426 6685 -1417
rect 6486 -1460 6493 -1426
rect 6673 -1460 6676 -1426
rect 6481 -1469 6493 -1460
rect 6545 -1469 6557 -1460
rect 6609 -1469 6621 -1460
rect 6673 -1469 6685 -1460
rect 6737 -1469 6749 -1417
rect 6801 -1469 6813 -1417
rect 6865 -1469 6877 -1417
rect 6929 -1426 6941 -1417
rect 6993 -1426 7005 -1417
rect 7057 -1426 7069 -1417
rect 7121 -1426 7133 -1417
rect 7185 -1426 7197 -1417
rect 6932 -1460 6941 -1426
rect 7185 -1460 7194 -1426
rect 6929 -1469 6941 -1460
rect 6993 -1469 7005 -1460
rect 7057 -1469 7069 -1460
rect 7121 -1469 7133 -1460
rect 7185 -1469 7197 -1460
rect 7249 -1469 7261 -1417
rect 7313 -1469 7325 -1417
rect 7377 -1469 7389 -1417
rect 7441 -1426 7453 -1417
rect 7505 -1426 7517 -1417
rect 7569 -1426 7581 -1417
rect 7633 -1426 7645 -1417
rect 7450 -1460 7453 -1426
rect 7633 -1460 7638 -1426
rect 7441 -1469 7453 -1460
rect 7505 -1469 7517 -1460
rect 7569 -1469 7581 -1460
rect 7633 -1469 7645 -1460
rect 7697 -1469 7709 -1417
rect 7761 -1469 7773 -1417
rect 7825 -1420 7831 -1417
rect 7825 -1466 7832 -1420
rect 7936 -1421 7942 -1387
rect 7976 -1421 7982 -1387
rect 7936 -1465 7982 -1421
rect 7825 -1469 7831 -1466
rect 5728 -1506 5734 -1472
rect 5768 -1506 5774 -1472
rect 5728 -1545 5774 -1506
rect 5728 -1579 5734 -1545
rect 5768 -1579 5774 -1545
rect 7936 -1499 7942 -1465
rect 7976 -1499 7982 -1465
rect 7936 -1543 7982 -1499
rect 5728 -1618 5774 -1579
rect 5728 -1652 5734 -1618
rect 5768 -1652 5774 -1618
rect 5840 -1625 5846 -1573
rect 5898 -1625 5911 -1573
rect 5963 -1625 5976 -1573
rect 6028 -1582 6041 -1573
rect 6093 -1582 6106 -1573
rect 6158 -1582 6171 -1573
rect 6223 -1582 6236 -1573
rect 6036 -1616 6041 -1582
rect 6223 -1616 6227 -1582
rect 6028 -1625 6041 -1616
rect 6093 -1625 6106 -1616
rect 6158 -1625 6171 -1616
rect 6223 -1625 6236 -1616
rect 6288 -1625 6301 -1573
rect 6353 -1625 6365 -1573
rect 6417 -1625 6429 -1573
rect 6481 -1582 6493 -1573
rect 6545 -1582 6557 -1573
rect 6609 -1582 6621 -1573
rect 6673 -1582 6685 -1573
rect 6486 -1616 6493 -1582
rect 6673 -1616 6676 -1582
rect 6481 -1625 6493 -1616
rect 6545 -1625 6557 -1616
rect 6609 -1625 6621 -1616
rect 6673 -1625 6685 -1616
rect 6737 -1625 6749 -1573
rect 6801 -1625 6813 -1573
rect 6865 -1625 6877 -1573
rect 6929 -1582 6941 -1573
rect 6993 -1582 7005 -1573
rect 7057 -1582 7069 -1573
rect 7121 -1582 7133 -1573
rect 7185 -1582 7197 -1573
rect 6932 -1616 6941 -1582
rect 7185 -1616 7194 -1582
rect 6929 -1625 6941 -1616
rect 6993 -1625 7005 -1616
rect 7057 -1625 7069 -1616
rect 7121 -1625 7133 -1616
rect 7185 -1625 7197 -1616
rect 7249 -1625 7261 -1573
rect 7313 -1625 7325 -1573
rect 7377 -1625 7389 -1573
rect 7441 -1582 7453 -1573
rect 7505 -1582 7517 -1573
rect 7569 -1582 7581 -1573
rect 7633 -1582 7645 -1573
rect 7450 -1616 7453 -1582
rect 7633 -1616 7638 -1582
rect 7441 -1625 7453 -1616
rect 7505 -1625 7517 -1616
rect 7569 -1625 7581 -1616
rect 7633 -1625 7645 -1616
rect 7697 -1625 7709 -1573
rect 7761 -1625 7773 -1573
rect 7825 -1576 7831 -1573
rect 7825 -1622 7832 -1576
rect 7936 -1577 7942 -1543
rect 7976 -1577 7982 -1543
rect 7936 -1622 7982 -1577
rect 7825 -1625 7831 -1622
rect 5728 -1691 5774 -1652
tri 7917 -1656 7936 -1637 se
rect 7936 -1656 7942 -1622
rect 7976 -1656 7982 -1622
rect 5728 -1725 5734 -1691
rect 5768 -1725 5774 -1691
rect 5728 -1764 5774 -1725
tri 7888 -1685 7917 -1656 se
rect 7917 -1685 7982 -1656
rect 7888 -1692 7982 -1685
rect 5728 -1798 5734 -1764
rect 5768 -1798 5774 -1764
rect 5840 -1781 5846 -1729
rect 5898 -1781 5911 -1729
rect 5963 -1781 5976 -1729
rect 6028 -1738 6041 -1729
rect 6093 -1738 6106 -1729
rect 6158 -1738 6171 -1729
rect 6223 -1738 6236 -1729
rect 6036 -1772 6041 -1738
rect 6223 -1772 6227 -1738
rect 6028 -1781 6041 -1772
rect 6093 -1781 6106 -1772
rect 6158 -1781 6171 -1772
rect 6223 -1781 6236 -1772
rect 6288 -1781 6301 -1729
rect 6353 -1781 6365 -1729
rect 6417 -1781 6429 -1729
rect 6481 -1738 6493 -1729
rect 6545 -1738 6557 -1729
rect 6609 -1738 6621 -1729
rect 6673 -1738 6685 -1729
rect 6486 -1772 6493 -1738
rect 6673 -1772 6676 -1738
rect 6481 -1781 6493 -1772
rect 6545 -1781 6557 -1772
rect 6609 -1781 6621 -1772
rect 6673 -1781 6685 -1772
rect 6737 -1781 6749 -1729
rect 6801 -1781 6813 -1729
rect 6865 -1781 6877 -1729
rect 6929 -1738 6941 -1729
rect 6993 -1738 7005 -1729
rect 7057 -1738 7069 -1729
rect 7121 -1738 7133 -1729
rect 7185 -1738 7197 -1729
rect 6932 -1772 6941 -1738
rect 7185 -1772 7194 -1738
rect 6929 -1781 6941 -1772
rect 6993 -1781 7005 -1772
rect 7057 -1781 7069 -1772
rect 7121 -1781 7133 -1772
rect 7185 -1781 7197 -1772
rect 7249 -1781 7261 -1729
rect 7313 -1781 7325 -1729
rect 7377 -1781 7389 -1729
rect 7441 -1738 7453 -1729
rect 7505 -1738 7517 -1729
rect 7569 -1738 7581 -1729
rect 7633 -1738 7645 -1729
rect 7450 -1772 7453 -1738
rect 7633 -1772 7638 -1738
rect 7441 -1781 7453 -1772
rect 7505 -1781 7517 -1772
rect 7569 -1781 7581 -1772
rect 7633 -1781 7645 -1772
rect 7697 -1781 7709 -1729
rect 7761 -1781 7773 -1729
rect 7825 -1732 7831 -1729
rect 7825 -1778 7832 -1732
rect 7888 -1744 7909 -1692
rect 7961 -1701 7982 -1692
rect 7976 -1735 7982 -1701
rect 7961 -1744 7982 -1735
rect 7888 -1766 7982 -1744
rect 7825 -1781 7831 -1778
rect 5728 -1837 5774 -1798
rect 5728 -1871 5734 -1837
rect 5768 -1871 5774 -1837
rect 5728 -1883 5774 -1871
rect 7888 -1818 7909 -1766
rect 7961 -1780 7982 -1766
rect 7976 -1814 7982 -1780
rect 7961 -1818 7982 -1814
rect 7888 -1841 7982 -1818
rect 5611 -1932 5657 -1888
rect 5611 -1966 5617 -1932
rect 5651 -1966 5657 -1932
rect 5840 -1937 5846 -1885
rect 5898 -1937 5911 -1885
rect 5963 -1937 5976 -1885
rect 6028 -1894 6041 -1885
rect 6093 -1894 6106 -1885
rect 6158 -1894 6171 -1885
rect 6223 -1894 6236 -1885
rect 6036 -1928 6041 -1894
rect 6223 -1928 6227 -1894
rect 6028 -1937 6041 -1928
rect 6093 -1937 6106 -1928
rect 6158 -1937 6171 -1928
rect 6223 -1937 6236 -1928
rect 6288 -1937 6301 -1885
rect 6353 -1937 6365 -1885
rect 6417 -1937 6429 -1885
rect 6481 -1894 6493 -1885
rect 6545 -1894 6557 -1885
rect 6609 -1894 6621 -1885
rect 6673 -1894 6685 -1885
rect 6486 -1928 6493 -1894
rect 6673 -1928 6676 -1894
rect 6481 -1937 6493 -1928
rect 6545 -1937 6557 -1928
rect 6609 -1937 6621 -1928
rect 6673 -1937 6685 -1928
rect 6737 -1937 6749 -1885
rect 6801 -1937 6813 -1885
rect 6865 -1937 6877 -1885
rect 6929 -1894 6941 -1885
rect 6993 -1894 7005 -1885
rect 7057 -1894 7069 -1885
rect 7121 -1894 7133 -1885
rect 7185 -1894 7197 -1885
rect 6932 -1928 6941 -1894
rect 7185 -1928 7194 -1894
rect 6929 -1937 6941 -1928
rect 6993 -1937 7005 -1928
rect 7057 -1937 7069 -1928
rect 7121 -1937 7133 -1928
rect 7185 -1937 7197 -1928
rect 7249 -1937 7261 -1885
rect 7313 -1937 7325 -1885
rect 7377 -1937 7389 -1885
rect 7441 -1894 7453 -1885
rect 7505 -1894 7517 -1885
rect 7569 -1894 7581 -1885
rect 7633 -1894 7645 -1885
rect 7450 -1928 7453 -1894
rect 7633 -1928 7638 -1894
rect 7441 -1937 7453 -1928
rect 7505 -1937 7517 -1928
rect 7569 -1937 7581 -1928
rect 7633 -1937 7645 -1928
rect 7697 -1937 7709 -1885
rect 7761 -1937 7773 -1885
rect 7825 -1888 7831 -1885
rect 7825 -1934 7832 -1888
rect 7888 -1893 7909 -1841
rect 7961 -1859 7982 -1841
rect 7976 -1893 7982 -1859
rect 7888 -1916 7982 -1893
rect 7825 -1937 7831 -1934
rect 5611 -2004 5657 -1966
rect 7888 -1968 7909 -1916
rect 7961 -1938 7982 -1916
rect 7888 -1972 7942 -1968
rect 7976 -1972 7982 -1938
tri 7862 -2004 7888 -1978 se
rect 7888 -1991 7982 -1972
rect 7888 -2004 7909 -1991
rect 5611 -2010 7909 -2004
rect 5611 -2044 5689 -2010
rect 5723 -2044 5762 -2010
rect 5796 -2044 5835 -2010
rect 5869 -2044 5908 -2010
rect 5942 -2044 5981 -2010
rect 6015 -2044 6054 -2010
rect 6088 -2044 6127 -2010
rect 6161 -2044 6200 -2010
rect 6234 -2044 6273 -2010
rect 6307 -2044 6346 -2010
rect 6380 -2044 6419 -2010
rect 6453 -2044 6492 -2010
rect 6526 -2044 6565 -2010
rect 6599 -2044 6638 -2010
rect 6672 -2044 6711 -2010
rect 6745 -2044 6784 -2010
rect 6818 -2044 6857 -2010
rect 6891 -2044 6930 -2010
rect 6964 -2044 7003 -2010
rect 7037 -2044 7076 -2010
rect 7110 -2044 7149 -2010
rect 7183 -2044 7222 -2010
rect 7256 -2044 7294 -2010
rect 7328 -2044 7366 -2010
rect 7400 -2044 7438 -2010
rect 7472 -2044 7510 -2010
rect 7544 -2044 7582 -2010
rect 7616 -2044 7654 -2010
rect 7688 -2044 7726 -2010
rect 7760 -2044 7798 -2010
rect 7832 -2044 7870 -2010
rect 7904 -2043 7909 -2010
rect 7961 -2043 7982 -1991
rect 7904 -2044 7982 -2043
rect 5611 -2050 7982 -2044
<< via1 >>
rect -358 1460 -322 1494
rect -322 1460 -306 1494
rect -294 1460 -288 1494
rect -288 1460 -242 1494
rect -358 1442 -306 1460
rect -294 1442 -242 1460
rect -358 1384 -306 1421
rect -294 1384 -242 1421
rect -358 1369 -322 1384
rect -322 1369 -306 1384
rect -294 1369 -288 1384
rect -288 1369 -242 1384
rect -358 1296 -306 1348
rect -294 1296 -242 1348
rect -490 851 -118 967
rect 320 935 324 967
rect 324 935 358 967
rect 358 935 396 967
rect 396 935 430 967
rect 430 935 436 967
rect 320 892 436 935
rect 320 858 324 892
rect 324 858 358 892
rect 358 858 396 892
rect 396 858 430 892
rect 430 858 436 892
rect 320 851 436 858
rect 640 1091 692 1143
rect 712 1091 764 1143
rect 784 1091 836 1143
rect 855 1091 907 1143
rect 640 1027 692 1079
rect 712 1027 764 1079
rect 784 1027 836 1079
rect 855 1027 907 1079
rect 1118 1081 1170 1133
rect 1195 1081 1247 1133
rect 1272 1081 1324 1133
rect 1348 1081 1400 1133
rect 1424 1081 1476 1133
rect 1500 1081 1552 1133
rect 1118 1042 1124 1055
rect 1124 1042 1158 1055
rect 1158 1042 1170 1055
rect 1118 1003 1170 1042
rect 1195 1042 1202 1055
rect 1202 1042 1236 1055
rect 1236 1042 1247 1055
rect 1195 1003 1247 1042
rect 1272 1042 1280 1055
rect 1280 1042 1314 1055
rect 1314 1042 1324 1055
rect 1272 1003 1324 1042
rect 1348 1042 1358 1055
rect 1358 1042 1392 1055
rect 1392 1042 1400 1055
rect 1348 1003 1400 1042
rect 1424 1042 1435 1055
rect 1435 1042 1469 1055
rect 1469 1042 1476 1055
rect 1424 1003 1476 1042
rect 1500 1042 1512 1055
rect 1512 1042 1546 1055
rect 1546 1042 1552 1055
rect 1500 1003 1552 1042
rect 640 790 692 796
rect 640 756 641 790
rect 641 756 675 790
rect 675 756 692 790
rect 640 744 692 756
rect 712 790 764 796
rect 712 756 716 790
rect 716 756 750 790
rect 750 756 764 790
rect 712 744 764 756
rect 784 790 836 796
rect 784 756 791 790
rect 791 756 825 790
rect 825 756 836 790
rect 784 744 836 756
rect 855 790 907 796
rect 855 756 866 790
rect 866 756 900 790
rect 900 756 907 790
rect 855 744 907 756
rect 467 594 519 598
rect 467 560 476 594
rect 476 560 510 594
rect 510 560 519 594
rect 467 546 519 560
rect 467 522 519 534
rect 467 488 476 522
rect 476 488 510 522
rect 510 488 519 522
rect 640 680 692 732
rect 712 680 764 732
rect 784 680 836 732
rect 855 680 907 732
rect 1117 634 1169 682
rect 1117 630 1123 634
rect 1123 630 1157 634
rect 1157 630 1169 634
rect 1194 634 1246 682
rect 1194 630 1201 634
rect 1201 630 1235 634
rect 1235 630 1246 634
rect 1271 634 1323 682
rect 1271 630 1279 634
rect 1279 630 1313 634
rect 1313 630 1323 634
rect 1348 634 1400 682
rect 1348 630 1357 634
rect 1357 630 1391 634
rect 1391 630 1400 634
rect 1424 634 1476 682
rect 1424 630 1435 634
rect 1435 630 1469 634
rect 1469 630 1476 634
rect 1500 634 1552 682
rect 1500 630 1512 634
rect 1512 630 1546 634
rect 1546 630 1552 634
rect 1117 600 1123 604
rect 1123 600 1157 604
rect 1157 600 1169 604
rect 1117 552 1169 600
rect 1194 600 1201 604
rect 1201 600 1235 604
rect 1235 600 1246 604
rect 1194 552 1246 600
rect 1271 600 1279 604
rect 1279 600 1313 604
rect 1313 600 1323 604
rect 1271 552 1323 600
rect 1348 600 1357 604
rect 1357 600 1391 604
rect 1391 600 1400 604
rect 1348 552 1400 600
rect 1424 600 1435 604
rect 1435 600 1469 604
rect 1469 600 1476 604
rect 1424 552 1476 600
rect 1500 600 1512 604
rect 1512 600 1546 604
rect 1546 600 1552 604
rect 1500 552 1552 600
rect 467 482 519 488
rect 3599 1450 3651 1456
rect 3665 1450 3717 1456
rect 3731 1450 3783 1456
rect 3797 1450 3849 1456
rect 3863 1450 3915 1456
rect 3929 1450 3981 1456
rect 3995 1450 4047 1456
rect 3599 1416 3624 1450
rect 3624 1416 3651 1450
rect 3665 1416 3697 1450
rect 3697 1416 3717 1450
rect 3731 1416 3770 1450
rect 3770 1416 3783 1450
rect 3797 1416 3804 1450
rect 3804 1416 3843 1450
rect 3843 1416 3849 1450
rect 3863 1416 3877 1450
rect 3877 1416 3915 1450
rect 3929 1416 3950 1450
rect 3950 1416 3981 1450
rect 3995 1416 4023 1450
rect 4023 1416 4047 1450
rect 3599 1404 3651 1416
rect 3665 1404 3717 1416
rect 3731 1404 3783 1416
rect 3797 1404 3849 1416
rect 3863 1404 3915 1416
rect 3929 1404 3981 1416
rect 3995 1404 4047 1416
rect 4061 1450 4113 1456
rect 4061 1416 4062 1450
rect 4062 1416 4096 1450
rect 4096 1416 4113 1450
rect 4061 1404 4113 1416
rect 4127 1450 4179 1456
rect 4127 1416 4135 1450
rect 4135 1416 4169 1450
rect 4169 1416 4179 1450
rect 4127 1404 4179 1416
rect 4193 1450 4245 1456
rect 4193 1416 4208 1450
rect 4208 1416 4242 1450
rect 4242 1416 4245 1450
rect 4193 1404 4245 1416
rect 4259 1450 4311 1456
rect 4325 1450 4377 1456
rect 4391 1450 4443 1456
rect 4457 1450 4509 1456
rect 4523 1450 4575 1456
rect 4589 1450 4641 1456
rect 4655 1450 4707 1456
rect 4721 1450 4773 1456
rect 4259 1416 4281 1450
rect 4281 1416 4311 1450
rect 4325 1416 4354 1450
rect 4354 1416 4377 1450
rect 4391 1416 4427 1450
rect 4427 1416 4443 1450
rect 4457 1416 4461 1450
rect 4461 1416 4500 1450
rect 4500 1416 4509 1450
rect 4523 1416 4534 1450
rect 4534 1416 4573 1450
rect 4573 1416 4575 1450
rect 4589 1416 4607 1450
rect 4607 1416 4641 1450
rect 4655 1416 4680 1450
rect 4680 1416 4707 1450
rect 4721 1416 4753 1450
rect 4753 1416 4773 1450
rect 4259 1404 4311 1416
rect 4325 1404 4377 1416
rect 4391 1404 4443 1416
rect 4457 1404 4509 1416
rect 4523 1404 4575 1416
rect 4589 1404 4641 1416
rect 4655 1404 4707 1416
rect 4721 1404 4773 1416
rect 4786 1450 4838 1456
rect 4786 1416 4792 1450
rect 4792 1416 4826 1450
rect 4826 1416 4838 1450
rect 4786 1404 4838 1416
rect 4851 1450 4903 1456
rect 4851 1416 4865 1450
rect 4865 1416 4899 1450
rect 4899 1416 4903 1450
rect 4851 1404 4903 1416
rect 4916 1450 4968 1456
rect 4981 1450 5033 1456
rect 5046 1450 5098 1456
rect 5111 1450 5163 1456
rect 5176 1450 5228 1456
rect 5241 1450 5293 1456
rect 4916 1416 4938 1450
rect 4938 1416 4968 1450
rect 4981 1416 5011 1450
rect 5011 1416 5033 1450
rect 5046 1416 5084 1450
rect 5084 1416 5098 1450
rect 5111 1416 5118 1450
rect 5118 1416 5157 1450
rect 5157 1416 5163 1450
rect 5176 1416 5191 1450
rect 5191 1416 5228 1450
rect 5241 1416 5264 1450
rect 5264 1416 5293 1450
rect 6644 1416 6661 1450
rect 6661 1416 6696 1450
rect 4916 1404 4968 1416
rect 4981 1404 5033 1416
rect 5046 1404 5098 1416
rect 5111 1404 5163 1416
rect 5176 1404 5228 1416
rect 5241 1404 5293 1416
rect 6644 1398 6696 1416
rect 6716 1398 6768 1450
rect 6788 1398 6840 1450
rect 3599 1378 3651 1392
rect 3665 1378 3717 1392
rect 3731 1378 3783 1392
rect 3797 1378 3849 1392
rect 3863 1378 3915 1392
rect 3929 1378 3981 1392
rect 3995 1378 4047 1392
rect 3599 1344 3624 1378
rect 3624 1344 3651 1378
rect 3665 1344 3697 1378
rect 3697 1344 3717 1378
rect 3731 1344 3770 1378
rect 3770 1344 3783 1378
rect 3797 1344 3804 1378
rect 3804 1344 3843 1378
rect 3843 1344 3849 1378
rect 3863 1344 3877 1378
rect 3877 1344 3915 1378
rect 3929 1344 3950 1378
rect 3950 1344 3981 1378
rect 3995 1344 4023 1378
rect 4023 1344 4047 1378
rect 3599 1340 3651 1344
rect 3665 1340 3717 1344
rect 3731 1340 3783 1344
rect 3797 1340 3849 1344
rect 3863 1340 3915 1344
rect 3929 1340 3981 1344
rect 3995 1340 4047 1344
rect 4061 1378 4113 1392
rect 4061 1344 4062 1378
rect 4062 1344 4096 1378
rect 4096 1344 4113 1378
rect 4061 1340 4113 1344
rect 4127 1378 4179 1392
rect 4127 1344 4135 1378
rect 4135 1344 4169 1378
rect 4169 1344 4179 1378
rect 4127 1340 4179 1344
rect 4193 1378 4245 1392
rect 4193 1344 4208 1378
rect 4208 1344 4242 1378
rect 4242 1344 4245 1378
rect 4193 1340 4245 1344
rect 4259 1378 4311 1392
rect 4325 1378 4377 1392
rect 4391 1378 4443 1392
rect 4457 1378 4509 1392
rect 4523 1378 4575 1392
rect 4589 1378 4641 1392
rect 4655 1378 4707 1392
rect 4721 1378 4773 1392
rect 4259 1344 4281 1378
rect 4281 1344 4311 1378
rect 4325 1344 4354 1378
rect 4354 1344 4377 1378
rect 4391 1344 4427 1378
rect 4427 1344 4443 1378
rect 4457 1344 4461 1378
rect 4461 1344 4500 1378
rect 4500 1344 4509 1378
rect 4523 1344 4534 1378
rect 4534 1344 4573 1378
rect 4573 1344 4575 1378
rect 4589 1344 4607 1378
rect 4607 1344 4641 1378
rect 4655 1344 4680 1378
rect 4680 1344 4707 1378
rect 4721 1344 4753 1378
rect 4753 1344 4773 1378
rect 4259 1340 4311 1344
rect 4325 1340 4377 1344
rect 4391 1340 4443 1344
rect 4457 1340 4509 1344
rect 4523 1340 4575 1344
rect 4589 1340 4641 1344
rect 4655 1340 4707 1344
rect 4721 1340 4773 1344
rect 4786 1378 4838 1392
rect 4786 1344 4792 1378
rect 4792 1344 4826 1378
rect 4826 1344 4838 1378
rect 4786 1340 4838 1344
rect 4851 1378 4903 1392
rect 4851 1344 4865 1378
rect 4865 1344 4899 1378
rect 4899 1344 4903 1378
rect 4851 1340 4903 1344
rect 4916 1378 4968 1392
rect 4981 1378 5033 1392
rect 5046 1378 5098 1392
rect 5111 1378 5163 1392
rect 5176 1378 5228 1392
rect 5241 1378 5293 1392
rect 6644 1378 6696 1379
rect 6716 1378 6768 1379
rect 4916 1344 4938 1378
rect 4938 1344 4968 1378
rect 4981 1344 5011 1378
rect 5011 1344 5033 1378
rect 5046 1344 5084 1378
rect 5084 1344 5098 1378
rect 5111 1344 5118 1378
rect 5118 1344 5157 1378
rect 5157 1344 5163 1378
rect 5176 1344 5191 1378
rect 5191 1344 5228 1378
rect 5241 1344 5264 1378
rect 5264 1344 5293 1378
rect 4916 1340 4968 1344
rect 4981 1340 5033 1344
rect 5046 1340 5098 1344
rect 5111 1340 5163 1344
rect 5176 1340 5228 1344
rect 5241 1340 5293 1344
rect 6644 1327 6696 1378
rect 6716 1327 6733 1378
rect 6733 1327 6768 1378
rect 6788 1327 6840 1379
rect 3136 1258 3188 1267
rect 3136 1224 3141 1258
rect 3141 1224 3175 1258
rect 3175 1224 3188 1258
rect 3136 1215 3188 1224
rect 3203 1258 3255 1267
rect 3203 1224 3215 1258
rect 3215 1224 3249 1258
rect 3249 1224 3255 1258
rect 3203 1215 3255 1224
rect 3269 1258 3321 1267
rect 3335 1258 3387 1267
rect 3401 1258 3453 1267
rect 3269 1224 3289 1258
rect 3289 1224 3321 1258
rect 3335 1224 3363 1258
rect 3363 1224 3387 1258
rect 3401 1224 3437 1258
rect 3437 1224 3453 1258
rect 3269 1215 3321 1224
rect 3335 1215 3387 1224
rect 3401 1215 3453 1224
rect 5820 1258 5872 1267
rect 5885 1258 5937 1267
rect 5949 1258 6001 1267
rect 5820 1224 5825 1258
rect 5825 1224 5865 1258
rect 5865 1224 5872 1258
rect 5885 1224 5899 1258
rect 5899 1224 5937 1258
rect 5949 1224 5973 1258
rect 5973 1224 6001 1258
rect 5820 1215 5872 1224
rect 5885 1215 5937 1224
rect 5949 1215 6001 1224
rect 6013 1258 6065 1267
rect 6013 1224 6047 1258
rect 6047 1224 6065 1258
rect 6013 1215 6065 1224
rect 6077 1258 6129 1267
rect 6077 1224 6087 1258
rect 6087 1224 6121 1258
rect 6121 1224 6129 1258
rect 6077 1215 6129 1224
rect 6141 1258 6193 1267
rect 6205 1258 6257 1267
rect 6269 1258 6321 1267
rect 6333 1258 6385 1267
rect 6397 1258 6449 1267
rect 6141 1224 6161 1258
rect 6161 1224 6193 1258
rect 6205 1224 6235 1258
rect 6235 1224 6257 1258
rect 6269 1224 6309 1258
rect 6309 1224 6321 1258
rect 6333 1224 6343 1258
rect 6343 1224 6383 1258
rect 6383 1224 6385 1258
rect 6397 1224 6417 1258
rect 6417 1224 6449 1258
rect 6141 1215 6193 1224
rect 6205 1215 6257 1224
rect 6269 1215 6321 1224
rect 6333 1215 6385 1224
rect 6397 1215 6449 1224
rect 2154 1125 2159 1141
rect 2159 1125 2193 1141
rect 2193 1125 2206 1141
rect 2154 1089 2206 1125
rect 2218 1125 2231 1141
rect 2231 1125 2265 1141
rect 2265 1125 2270 1141
rect 2218 1089 2270 1125
rect 2154 1052 2159 1075
rect 2159 1052 2193 1075
rect 2193 1052 2206 1075
rect 2154 1023 2206 1052
rect 2218 1052 2231 1075
rect 2231 1052 2265 1075
rect 2265 1052 2270 1075
rect 2218 1023 2270 1052
rect 2154 979 2159 1009
rect 2159 979 2193 1009
rect 2193 979 2206 1009
rect 2154 957 2206 979
rect 2218 979 2231 1009
rect 2231 979 2265 1009
rect 2265 979 2270 1009
rect 2218 957 2270 979
rect 2305 1201 2357 1207
rect 2305 1167 2311 1201
rect 2311 1167 2345 1201
rect 2345 1167 2357 1201
rect 2305 1155 2357 1167
rect 2305 1128 2357 1134
rect 6539 1212 6591 1264
rect 6539 1167 6547 1191
rect 6547 1167 6581 1191
rect 6581 1167 6591 1191
rect 6539 1139 6591 1167
rect 2305 1094 2311 1128
rect 2311 1094 2345 1128
rect 2345 1094 2357 1128
rect 2305 1082 2357 1094
rect 3599 1102 3651 1111
rect 3670 1102 3722 1111
rect 3741 1102 3793 1111
rect 3811 1102 3863 1111
rect 3881 1102 3933 1111
rect 3951 1102 4003 1111
rect 3599 1068 3617 1102
rect 3617 1068 3651 1102
rect 3670 1068 3690 1102
rect 3690 1068 3722 1102
rect 3741 1068 3763 1102
rect 3763 1068 3793 1102
rect 3811 1068 3836 1102
rect 3836 1068 3863 1102
rect 3881 1068 3909 1102
rect 3909 1068 3933 1102
rect 3951 1068 3982 1102
rect 3982 1068 4003 1102
rect 2305 1055 2357 1061
rect 3599 1059 3651 1068
rect 3670 1059 3722 1068
rect 3741 1059 3793 1068
rect 3811 1059 3863 1068
rect 3881 1059 3933 1068
rect 3951 1059 4003 1068
rect 4021 1102 4073 1111
rect 4021 1068 4055 1102
rect 4055 1068 4073 1102
rect 4021 1059 4073 1068
rect 4091 1102 4143 1111
rect 4091 1068 4094 1102
rect 4094 1068 4128 1102
rect 4128 1068 4143 1102
rect 4091 1059 4143 1068
rect 4161 1102 4213 1111
rect 4161 1068 4167 1102
rect 4167 1068 4201 1102
rect 4201 1068 4213 1102
rect 4161 1059 4213 1068
rect 4231 1102 4283 1111
rect 4231 1068 4240 1102
rect 4240 1068 4274 1102
rect 4274 1068 4283 1102
rect 4231 1059 4283 1068
rect 4301 1102 4353 1111
rect 4301 1068 4313 1102
rect 4313 1068 4347 1102
rect 4347 1068 4353 1102
rect 4301 1059 4353 1068
rect 4539 1102 4591 1111
rect 4539 1068 4545 1102
rect 4545 1068 4579 1102
rect 4579 1068 4591 1102
rect 4539 1059 4591 1068
rect 4609 1102 4661 1111
rect 4609 1068 4618 1102
rect 4618 1068 4652 1102
rect 4652 1068 4661 1102
rect 4609 1059 4661 1068
rect 4679 1102 4731 1111
rect 4679 1068 4691 1102
rect 4691 1068 4725 1102
rect 4725 1068 4731 1102
rect 4679 1059 4731 1068
rect 4749 1102 4801 1111
rect 4749 1068 4764 1102
rect 4764 1068 4798 1102
rect 4798 1068 4801 1102
rect 4749 1059 4801 1068
rect 4819 1102 4871 1111
rect 4819 1068 4837 1102
rect 4837 1068 4871 1102
rect 4819 1059 4871 1068
rect 4889 1102 4941 1111
rect 4959 1102 5011 1111
rect 5029 1102 5081 1111
rect 5099 1102 5151 1111
rect 5170 1102 5222 1111
rect 5241 1102 5293 1111
rect 6162 1102 6214 1111
rect 6250 1102 6302 1111
rect 6338 1102 6390 1111
rect 4889 1068 4910 1102
rect 4910 1068 4941 1102
rect 4959 1068 4983 1102
rect 4983 1068 5011 1102
rect 5029 1068 5056 1102
rect 5056 1068 5081 1102
rect 5099 1068 5129 1102
rect 5129 1068 5151 1102
rect 5170 1068 5202 1102
rect 5202 1068 5222 1102
rect 5241 1068 5275 1102
rect 5275 1068 5293 1102
rect 6162 1068 6195 1102
rect 6195 1068 6214 1102
rect 6250 1068 6269 1102
rect 6269 1068 6302 1102
rect 6338 1068 6343 1102
rect 6343 1068 6383 1102
rect 6383 1068 6390 1102
rect 4889 1059 4941 1068
rect 4959 1059 5011 1068
rect 5029 1059 5081 1068
rect 5099 1059 5151 1068
rect 5170 1059 5222 1068
rect 5241 1059 5293 1068
rect 6162 1059 6214 1068
rect 6250 1059 6302 1068
rect 6338 1059 6390 1068
rect 2305 1021 2311 1055
rect 2311 1021 2345 1055
rect 2345 1021 2357 1055
rect 2305 1009 2357 1021
rect 2305 981 2357 988
rect 2305 947 2311 981
rect 2311 947 2345 981
rect 2345 947 2357 981
rect 2305 936 2357 947
rect 2305 907 2357 915
rect 2305 873 2311 907
rect 2311 873 2345 907
rect 2345 873 2357 907
rect 3136 946 3188 955
rect 3136 912 3141 946
rect 3141 912 3175 946
rect 3175 912 3188 946
rect 3136 903 3188 912
rect 3203 946 3255 955
rect 3203 912 3215 946
rect 3215 912 3249 946
rect 3249 912 3255 946
rect 3203 903 3255 912
rect 3269 946 3321 955
rect 3335 946 3387 955
rect 3401 946 3453 955
rect 3269 912 3289 946
rect 3289 912 3321 946
rect 3335 912 3363 946
rect 3363 912 3387 946
rect 3401 912 3437 946
rect 3437 912 3453 946
rect 3269 903 3321 912
rect 3335 903 3387 912
rect 3401 903 3453 912
rect 5820 946 5872 955
rect 5885 946 5937 955
rect 5949 946 6001 955
rect 5820 912 5825 946
rect 5825 912 5865 946
rect 5865 912 5872 946
rect 5885 912 5899 946
rect 5899 912 5937 946
rect 5949 912 5973 946
rect 5973 912 6001 946
rect 5820 903 5872 912
rect 5885 903 5937 912
rect 5949 903 6001 912
rect 6013 946 6065 955
rect 6013 912 6047 946
rect 6047 912 6065 946
rect 6013 903 6065 912
rect 6077 946 6129 955
rect 6077 912 6087 946
rect 6087 912 6121 946
rect 6121 912 6129 946
rect 6077 903 6129 912
rect 6141 946 6193 955
rect 6205 946 6257 955
rect 6269 946 6321 955
rect 6333 946 6385 955
rect 6397 946 6449 955
rect 6141 912 6161 946
rect 6161 912 6193 946
rect 6205 912 6235 946
rect 6235 912 6257 946
rect 6269 912 6309 946
rect 6309 912 6321 946
rect 6333 912 6343 946
rect 6343 912 6383 946
rect 6383 912 6385 946
rect 6397 912 6417 946
rect 6417 912 6449 946
rect 6141 903 6193 912
rect 6205 903 6257 912
rect 6269 903 6321 912
rect 6333 903 6385 912
rect 6397 903 6449 912
rect 2305 863 2357 873
rect 2305 833 2357 842
rect 2305 799 2311 833
rect 2311 799 2345 833
rect 2345 799 2357 833
rect 2305 790 2357 799
rect 2305 759 2357 769
rect 2305 725 2311 759
rect 2311 725 2345 759
rect 2345 725 2357 759
rect 3599 790 3651 799
rect 3670 790 3722 799
rect 3741 790 3793 799
rect 3811 790 3863 799
rect 3881 790 3933 799
rect 3951 790 4003 799
rect 3599 756 3617 790
rect 3617 756 3651 790
rect 3670 756 3690 790
rect 3690 756 3722 790
rect 3741 756 3763 790
rect 3763 756 3793 790
rect 3811 756 3836 790
rect 3836 756 3863 790
rect 3881 756 3909 790
rect 3909 756 3933 790
rect 3951 756 3982 790
rect 3982 756 4003 790
rect 3599 747 3651 756
rect 3670 747 3722 756
rect 3741 747 3793 756
rect 3811 747 3863 756
rect 3881 747 3933 756
rect 3951 747 4003 756
rect 4021 790 4073 799
rect 4021 756 4055 790
rect 4055 756 4073 790
rect 4021 747 4073 756
rect 4091 790 4143 799
rect 4091 756 4094 790
rect 4094 756 4128 790
rect 4128 756 4143 790
rect 4091 747 4143 756
rect 4161 790 4213 799
rect 4161 756 4167 790
rect 4167 756 4201 790
rect 4201 756 4213 790
rect 4161 747 4213 756
rect 4231 790 4283 799
rect 4231 756 4240 790
rect 4240 756 4274 790
rect 4274 756 4283 790
rect 4231 747 4283 756
rect 4301 790 4353 799
rect 4301 756 4313 790
rect 4313 756 4347 790
rect 4347 756 4353 790
rect 4301 747 4353 756
rect 4539 790 4591 799
rect 4539 756 4545 790
rect 4545 756 4579 790
rect 4579 756 4591 790
rect 4539 747 4591 756
rect 4609 790 4661 799
rect 4609 756 4618 790
rect 4618 756 4652 790
rect 4652 756 4661 790
rect 4609 747 4661 756
rect 4679 790 4731 799
rect 4679 756 4691 790
rect 4691 756 4725 790
rect 4725 756 4731 790
rect 4679 747 4731 756
rect 4749 790 4801 799
rect 4749 756 4764 790
rect 4764 756 4798 790
rect 4798 756 4801 790
rect 4749 747 4801 756
rect 4819 790 4871 799
rect 4819 756 4837 790
rect 4837 756 4871 790
rect 4819 747 4871 756
rect 4889 790 4941 799
rect 4959 790 5011 799
rect 5029 790 5081 799
rect 5099 790 5151 799
rect 5170 790 5222 799
rect 5241 790 5293 799
rect 6162 790 6214 799
rect 6250 790 6302 799
rect 6338 790 6390 799
rect 4889 756 4910 790
rect 4910 756 4941 790
rect 4959 756 4983 790
rect 4983 756 5011 790
rect 5029 756 5056 790
rect 5056 756 5081 790
rect 5099 756 5129 790
rect 5129 756 5151 790
rect 5170 756 5202 790
rect 5202 756 5222 790
rect 5241 756 5275 790
rect 5275 756 5293 790
rect 6162 756 6195 790
rect 6195 756 6214 790
rect 6250 756 6269 790
rect 6269 756 6302 790
rect 6338 756 6343 790
rect 6343 756 6383 790
rect 6383 756 6390 790
rect 4889 747 4941 756
rect 4959 747 5011 756
rect 5029 747 5081 756
rect 5099 747 5151 756
rect 5170 747 5222 756
rect 5241 747 5293 756
rect 6162 747 6214 756
rect 6250 747 6302 756
rect 6338 747 6390 756
rect 2305 717 2357 725
rect 2305 685 2357 697
rect 2305 651 2311 685
rect 2311 651 2345 685
rect 2345 651 2357 685
rect 2305 645 2357 651
rect 6539 691 6591 704
rect 6539 657 6547 691
rect 6547 657 6581 691
rect 6581 657 6591 691
rect 6539 652 6591 657
rect 3136 634 3188 643
rect 3136 600 3141 634
rect 3141 600 3175 634
rect 3175 600 3188 634
rect 3136 591 3188 600
rect 3203 634 3255 643
rect 3203 600 3215 634
rect 3215 600 3249 634
rect 3249 600 3255 634
rect 3203 591 3255 600
rect 3269 634 3321 643
rect 3335 634 3387 643
rect 3401 634 3453 643
rect 3269 600 3289 634
rect 3289 600 3321 634
rect 3335 600 3363 634
rect 3363 600 3387 634
rect 3401 600 3437 634
rect 3437 600 3453 634
rect 3269 591 3321 600
rect 3335 591 3387 600
rect 3401 591 3453 600
rect 5820 634 5872 643
rect 5885 634 5937 643
rect 5949 634 6001 643
rect 5820 600 5825 634
rect 5825 600 5865 634
rect 5865 600 5872 634
rect 5885 600 5899 634
rect 5899 600 5937 634
rect 5949 600 5973 634
rect 5973 600 6001 634
rect 5820 591 5872 600
rect 5885 591 5937 600
rect 5949 591 6001 600
rect 6013 634 6065 643
rect 6013 600 6047 634
rect 6047 600 6065 634
rect 6013 591 6065 600
rect 6077 634 6129 643
rect 6077 600 6087 634
rect 6087 600 6121 634
rect 6121 600 6129 634
rect 6077 591 6129 600
rect 6141 634 6193 643
rect 6205 634 6257 643
rect 6269 634 6321 643
rect 6333 634 6385 643
rect 6397 634 6449 643
rect 6141 600 6161 634
rect 6161 600 6193 634
rect 6205 600 6235 634
rect 6235 600 6257 634
rect 6269 600 6309 634
rect 6309 600 6321 634
rect 6333 600 6343 634
rect 6343 600 6383 634
rect 6383 600 6385 634
rect 6397 600 6417 634
rect 6417 600 6449 634
rect 6141 591 6193 600
rect 6205 591 6257 600
rect 6269 591 6321 600
rect 6333 591 6385 600
rect 6397 591 6449 600
rect 6539 579 6591 631
rect 3599 478 3651 487
rect 3670 478 3722 487
rect 3741 478 3793 487
rect 3811 478 3863 487
rect 3881 478 3933 487
rect 3951 478 4003 487
rect 3599 444 3617 478
rect 3617 444 3651 478
rect 3670 444 3690 478
rect 3690 444 3722 478
rect 3741 444 3763 478
rect 3763 444 3793 478
rect 3811 444 3836 478
rect 3836 444 3863 478
rect 3881 444 3909 478
rect 3909 444 3933 478
rect 3951 444 3982 478
rect 3982 444 4003 478
rect 3599 435 3651 444
rect 3670 435 3722 444
rect 3741 435 3793 444
rect 3811 435 3863 444
rect 3881 435 3933 444
rect 3951 435 4003 444
rect 4021 478 4073 487
rect 4021 444 4055 478
rect 4055 444 4073 478
rect 4021 435 4073 444
rect 4091 478 4143 487
rect 4091 444 4094 478
rect 4094 444 4128 478
rect 4128 444 4143 478
rect 4091 435 4143 444
rect 4161 478 4213 487
rect 4161 444 4167 478
rect 4167 444 4201 478
rect 4201 444 4213 478
rect 4161 435 4213 444
rect 4231 478 4283 487
rect 4231 444 4240 478
rect 4240 444 4274 478
rect 4274 444 4283 478
rect 4231 435 4283 444
rect 4301 478 4353 487
rect 4301 444 4313 478
rect 4313 444 4347 478
rect 4347 444 4353 478
rect 4301 435 4353 444
rect 4539 478 4591 487
rect 4539 444 4545 478
rect 4545 444 4579 478
rect 4579 444 4591 478
rect 4539 435 4591 444
rect 4609 478 4661 487
rect 4609 444 4618 478
rect 4618 444 4652 478
rect 4652 444 4661 478
rect 4609 435 4661 444
rect 4679 478 4731 487
rect 4679 444 4691 478
rect 4691 444 4725 478
rect 4725 444 4731 478
rect 4679 435 4731 444
rect 4749 478 4801 487
rect 4749 444 4764 478
rect 4764 444 4798 478
rect 4798 444 4801 478
rect 4749 435 4801 444
rect 4819 478 4871 487
rect 4819 444 4837 478
rect 4837 444 4871 478
rect 4819 435 4871 444
rect 4889 478 4941 487
rect 4959 478 5011 487
rect 5029 478 5081 487
rect 5099 478 5151 487
rect 5170 478 5222 487
rect 5241 478 5293 487
rect 4889 444 4910 478
rect 4910 444 4941 478
rect 4959 444 4983 478
rect 4983 444 5011 478
rect 5029 444 5056 478
rect 5056 444 5081 478
rect 5099 444 5129 478
rect 5129 444 5151 478
rect 5170 444 5202 478
rect 5202 444 5222 478
rect 5241 444 5275 478
rect 5275 444 5293 478
rect 6183 444 6195 456
rect 6195 444 6235 456
rect 6235 444 6269 456
rect 6269 444 6309 456
rect 6309 444 6343 456
rect 6343 444 6363 456
rect 4889 435 4941 444
rect 4959 435 5011 444
rect 5029 435 5081 444
rect 5099 435 5151 444
rect 5170 435 5222 444
rect 5241 435 5293 444
rect 3599 362 3651 414
rect 3665 362 3717 414
rect 3731 362 3783 414
rect 3797 362 3849 414
rect 3863 362 3915 414
rect 3929 362 3981 414
rect 3995 362 4047 414
rect 4061 362 4113 414
rect 4127 362 4179 414
rect 4193 362 4245 414
rect 4259 362 4311 414
rect 4325 362 4377 414
rect 4391 362 4443 414
rect 4457 362 4509 414
rect 4523 362 4575 414
rect 4589 362 4641 414
rect 4655 362 4707 414
rect 4721 362 4773 414
rect 4786 362 4838 414
rect 4851 362 4903 414
rect 4916 362 4968 414
rect 4981 362 5033 414
rect 5046 362 5098 414
rect 5111 362 5163 414
rect 5176 362 5228 414
rect 5241 362 5293 414
rect 6183 358 6363 444
rect 6183 340 6363 358
rect 8618 1450 8670 1456
rect 8684 1450 8736 1456
rect 8750 1450 8802 1456
rect 8816 1450 8868 1456
rect 8882 1450 8934 1456
rect 8948 1450 9000 1456
rect 9014 1450 9066 1456
rect 9080 1450 9132 1456
rect 9146 1450 9198 1456
rect 9212 1450 9264 1456
rect 9278 1450 9330 1456
rect 9344 1450 9396 1456
rect 9410 1450 9462 1456
rect 9476 1450 9528 1456
rect 9542 1450 9594 1456
rect 9608 1450 9660 1456
rect 9674 1450 9726 1456
rect 9740 1450 9792 1456
rect 9805 1450 9857 1456
rect 9870 1450 9922 1456
rect 9935 1450 9987 1456
rect 10000 1450 10052 1456
rect 10065 1450 10117 1456
rect 10130 1450 10182 1456
rect 10195 1450 10247 1456
rect 10260 1450 10312 1456
rect 8618 1404 8670 1450
rect 8684 1404 8736 1450
rect 8750 1404 8802 1450
rect 8816 1404 8868 1450
rect 8882 1404 8934 1450
rect 8948 1404 9000 1450
rect 9014 1404 9066 1450
rect 9080 1404 9132 1450
rect 9146 1404 9198 1450
rect 9212 1404 9264 1450
rect 9278 1404 9330 1450
rect 9344 1404 9396 1450
rect 9410 1404 9462 1450
rect 9476 1404 9528 1450
rect 9542 1404 9594 1450
rect 9608 1404 9660 1450
rect 9674 1404 9726 1450
rect 9740 1404 9792 1450
rect 9805 1404 9857 1450
rect 9870 1404 9922 1450
rect 9935 1404 9987 1450
rect 10000 1404 10052 1450
rect 10065 1404 10117 1450
rect 10130 1404 10182 1450
rect 10195 1404 10247 1450
rect 10260 1404 10312 1450
rect 8618 1344 8670 1392
rect 8684 1344 8736 1392
rect 8750 1344 8802 1392
rect 8816 1344 8868 1392
rect 8882 1344 8934 1392
rect 8948 1344 9000 1392
rect 9014 1344 9066 1392
rect 9080 1344 9132 1392
rect 9146 1344 9198 1392
rect 9212 1344 9264 1392
rect 9278 1344 9330 1392
rect 9344 1344 9396 1392
rect 9410 1344 9462 1392
rect 9476 1344 9528 1392
rect 9542 1344 9594 1392
rect 9608 1344 9660 1392
rect 9674 1344 9726 1392
rect 9740 1344 9792 1392
rect 9805 1344 9857 1392
rect 9870 1344 9922 1392
rect 9935 1344 9987 1392
rect 10000 1344 10052 1392
rect 10065 1344 10117 1392
rect 10130 1344 10182 1392
rect 10195 1344 10247 1392
rect 10260 1344 10312 1392
rect 8618 1340 8670 1344
rect 8684 1340 8736 1344
rect 8750 1340 8802 1344
rect 8816 1340 8868 1344
rect 8882 1340 8934 1344
rect 8948 1340 9000 1344
rect 9014 1340 9066 1344
rect 9080 1340 9132 1344
rect 9146 1340 9198 1344
rect 9212 1340 9264 1344
rect 9278 1340 9330 1344
rect 9344 1340 9396 1344
rect 9410 1340 9462 1344
rect 9476 1340 9528 1344
rect 9542 1340 9594 1344
rect 9608 1340 9660 1344
rect 9674 1340 9726 1344
rect 9740 1340 9792 1344
rect 9805 1340 9857 1344
rect 9870 1340 9922 1344
rect 9935 1340 9987 1344
rect 10000 1340 10052 1344
rect 10065 1340 10117 1344
rect 10130 1340 10182 1344
rect 10195 1340 10247 1344
rect 10260 1340 10312 1344
rect 7424 1258 7476 1267
rect 7496 1258 7548 1267
rect 7424 1224 7454 1258
rect 7454 1224 7476 1258
rect 7496 1224 7528 1258
rect 7528 1224 7548 1258
rect 7424 1215 7476 1224
rect 7496 1215 7548 1224
rect 7568 1258 7620 1267
rect 7568 1224 7602 1258
rect 7602 1224 7620 1258
rect 7568 1215 7620 1224
rect 7639 1258 7691 1267
rect 7639 1224 7642 1258
rect 7642 1224 7676 1258
rect 7676 1224 7691 1258
rect 7639 1215 7691 1224
rect 7710 1258 7762 1267
rect 7710 1224 7716 1258
rect 7716 1224 7750 1258
rect 7750 1224 7762 1258
rect 7710 1215 7762 1224
rect 7781 1258 7833 1267
rect 7781 1224 7790 1258
rect 7790 1224 7824 1258
rect 7824 1224 7833 1258
rect 7781 1215 7833 1224
rect 7852 1258 7904 1267
rect 7852 1224 7864 1258
rect 7864 1224 7898 1258
rect 7898 1224 7904 1258
rect 7852 1215 7904 1224
rect 7923 1258 7975 1267
rect 7923 1224 7938 1258
rect 7938 1224 7972 1258
rect 7972 1224 7975 1258
rect 7923 1215 7975 1224
rect 7994 1258 8046 1267
rect 7994 1224 8012 1258
rect 8012 1224 8046 1258
rect 7994 1215 8046 1224
rect 10458 1258 10510 1267
rect 10525 1258 10577 1267
rect 10591 1258 10643 1267
rect 10458 1224 10474 1258
rect 10474 1224 10510 1258
rect 10525 1224 10548 1258
rect 10548 1224 10577 1258
rect 10591 1224 10622 1258
rect 10622 1224 10643 1258
rect 10458 1215 10510 1224
rect 10525 1215 10577 1224
rect 10591 1215 10643 1224
rect 10657 1258 10709 1267
rect 10657 1224 10662 1258
rect 10662 1224 10696 1258
rect 10696 1224 10709 1258
rect 10657 1215 10709 1224
rect 10723 1258 10775 1267
rect 10723 1224 10736 1258
rect 10736 1224 10770 1258
rect 10770 1224 10775 1258
rect 10723 1215 10775 1224
rect 7322 1201 7374 1207
rect 7322 1167 7330 1201
rect 7330 1167 7364 1201
rect 7364 1167 7374 1201
rect 7322 1155 7374 1167
rect 7322 1127 7374 1141
rect 7322 1093 7330 1127
rect 7330 1093 7364 1127
rect 7364 1093 7374 1127
rect 11558 1201 11610 1207
rect 11558 1167 11566 1201
rect 11566 1167 11600 1201
rect 11600 1167 11610 1201
rect 11558 1155 11610 1167
rect 11558 1127 11610 1141
rect 7322 1089 7374 1093
rect 7322 1053 7374 1075
rect 8618 1102 8670 1111
rect 8689 1102 8741 1111
rect 8760 1102 8812 1111
rect 8830 1102 8882 1111
rect 8900 1102 8952 1111
rect 8970 1102 9022 1111
rect 8618 1068 8636 1102
rect 8636 1068 8670 1102
rect 8689 1068 8709 1102
rect 8709 1068 8741 1102
rect 8760 1068 8782 1102
rect 8782 1068 8812 1102
rect 8830 1068 8855 1102
rect 8855 1068 8882 1102
rect 8900 1068 8928 1102
rect 8928 1068 8952 1102
rect 8970 1068 9001 1102
rect 9001 1068 9022 1102
rect 8618 1059 8670 1068
rect 8689 1059 8741 1068
rect 8760 1059 8812 1068
rect 8830 1059 8882 1068
rect 8900 1059 8952 1068
rect 8970 1059 9022 1068
rect 9040 1102 9092 1111
rect 9040 1068 9074 1102
rect 9074 1068 9092 1102
rect 9040 1059 9092 1068
rect 9110 1102 9162 1111
rect 9110 1068 9113 1102
rect 9113 1068 9147 1102
rect 9147 1068 9162 1102
rect 9110 1059 9162 1068
rect 9180 1102 9232 1111
rect 9180 1068 9186 1102
rect 9186 1068 9220 1102
rect 9220 1068 9232 1102
rect 9180 1059 9232 1068
rect 9250 1102 9302 1111
rect 9250 1068 9259 1102
rect 9259 1068 9293 1102
rect 9293 1068 9302 1102
rect 9250 1059 9302 1068
rect 9320 1102 9372 1111
rect 9320 1068 9332 1102
rect 9332 1068 9366 1102
rect 9366 1068 9372 1102
rect 9320 1059 9372 1068
rect 9558 1102 9610 1111
rect 9558 1068 9564 1102
rect 9564 1068 9598 1102
rect 9598 1068 9610 1102
rect 9558 1059 9610 1068
rect 9628 1102 9680 1111
rect 9628 1068 9637 1102
rect 9637 1068 9671 1102
rect 9671 1068 9680 1102
rect 9628 1059 9680 1068
rect 9698 1102 9750 1111
rect 9698 1068 9710 1102
rect 9710 1068 9744 1102
rect 9744 1068 9750 1102
rect 9698 1059 9750 1068
rect 9768 1102 9820 1111
rect 9768 1068 9783 1102
rect 9783 1068 9817 1102
rect 9817 1068 9820 1102
rect 9768 1059 9820 1068
rect 9838 1102 9890 1111
rect 9838 1068 9856 1102
rect 9856 1068 9890 1102
rect 9838 1059 9890 1068
rect 9908 1102 9960 1111
rect 9978 1102 10030 1111
rect 10048 1102 10100 1111
rect 10118 1102 10170 1111
rect 10189 1102 10241 1111
rect 10260 1102 10312 1111
rect 9908 1068 9929 1102
rect 9929 1068 9960 1102
rect 9978 1068 10002 1102
rect 10002 1068 10030 1102
rect 10048 1068 10075 1102
rect 10075 1068 10100 1102
rect 10118 1068 10148 1102
rect 10148 1068 10170 1102
rect 10189 1068 10221 1102
rect 10221 1068 10241 1102
rect 10260 1068 10294 1102
rect 10294 1068 10312 1102
rect 9908 1059 9960 1068
rect 9978 1059 10030 1068
rect 10048 1059 10100 1068
rect 10118 1059 10170 1068
rect 10189 1059 10241 1068
rect 10260 1059 10312 1068
rect 11558 1093 11566 1127
rect 11566 1093 11600 1127
rect 11600 1093 11610 1127
rect 11558 1089 11610 1093
rect 7322 1023 7330 1053
rect 7330 1023 7364 1053
rect 7364 1023 7374 1053
rect 7322 979 7374 1009
rect 7322 957 7330 979
rect 7330 957 7364 979
rect 7364 957 7374 979
rect 11558 1053 11610 1075
rect 11558 1023 11566 1053
rect 11566 1023 11600 1053
rect 11600 1023 11610 1053
rect 11558 979 11610 1009
rect 11558 957 11566 979
rect 11566 957 11600 979
rect 11600 957 11610 979
rect 7322 905 7374 943
rect 7424 946 7476 955
rect 7495 946 7547 955
rect 7424 912 7454 946
rect 7454 912 7476 946
rect 7495 912 7528 946
rect 7528 912 7547 946
rect 7322 891 7330 905
rect 7330 891 7364 905
rect 7364 891 7374 905
rect 7424 903 7476 912
rect 7495 903 7547 912
rect 7566 946 7618 955
rect 7566 912 7568 946
rect 7568 912 7602 946
rect 7602 912 7618 946
rect 7566 903 7618 912
rect 7637 946 7689 955
rect 7637 912 7642 946
rect 7642 912 7676 946
rect 7676 912 7689 946
rect 7637 903 7689 912
rect 7707 946 7759 955
rect 7707 912 7716 946
rect 7716 912 7750 946
rect 7750 912 7759 946
rect 7707 903 7759 912
rect 7777 946 7829 955
rect 7777 912 7790 946
rect 7790 912 7824 946
rect 7824 912 7829 946
rect 7777 903 7829 912
rect 7847 946 7899 955
rect 7847 912 7864 946
rect 7864 912 7898 946
rect 7898 912 7899 946
rect 7847 903 7899 912
rect 7917 946 7969 955
rect 7987 946 8039 955
rect 7917 912 7938 946
rect 7938 912 7969 946
rect 7987 912 8012 946
rect 8012 912 8039 946
rect 7917 903 7969 912
rect 7987 903 8039 912
rect 10458 946 10510 955
rect 10525 946 10577 955
rect 10591 946 10643 955
rect 10458 912 10474 946
rect 10474 912 10510 946
rect 10525 912 10548 946
rect 10548 912 10577 946
rect 10591 912 10622 946
rect 10622 912 10643 946
rect 10458 903 10510 912
rect 10525 903 10577 912
rect 10591 903 10643 912
rect 10657 946 10709 955
rect 10657 912 10662 946
rect 10662 912 10696 946
rect 10696 912 10709 946
rect 10657 903 10709 912
rect 10723 946 10775 955
rect 10723 912 10736 946
rect 10736 912 10770 946
rect 10770 912 10775 946
rect 10723 903 10775 912
rect 11558 905 11610 943
rect 7322 871 7330 877
rect 7330 871 7364 877
rect 7364 871 7374 877
rect 7322 831 7374 871
rect 7322 825 7330 831
rect 7330 825 7364 831
rect 7364 825 7374 831
rect 7322 797 7330 811
rect 7330 797 7364 811
rect 7364 797 7374 811
rect 11558 891 11566 905
rect 11566 891 11600 905
rect 11600 891 11610 905
rect 11558 871 11566 877
rect 11566 871 11600 877
rect 11600 871 11610 877
rect 11558 831 11610 871
rect 11558 825 11566 831
rect 11566 825 11600 831
rect 11600 825 11610 831
rect 7322 759 7374 797
rect 8618 790 8670 799
rect 8689 790 8741 799
rect 8760 790 8812 799
rect 8830 790 8882 799
rect 8900 790 8952 799
rect 8970 790 9022 799
rect 8618 756 8636 790
rect 8636 756 8670 790
rect 8689 756 8709 790
rect 8709 756 8741 790
rect 8760 756 8782 790
rect 8782 756 8812 790
rect 8830 756 8855 790
rect 8855 756 8882 790
rect 8900 756 8928 790
rect 8928 756 8952 790
rect 8970 756 9001 790
rect 9001 756 9022 790
rect 8618 747 8670 756
rect 8689 747 8741 756
rect 8760 747 8812 756
rect 8830 747 8882 756
rect 8900 747 8952 756
rect 8970 747 9022 756
rect 9040 790 9092 799
rect 9040 756 9074 790
rect 9074 756 9092 790
rect 9040 747 9092 756
rect 9110 790 9162 799
rect 9110 756 9113 790
rect 9113 756 9147 790
rect 9147 756 9162 790
rect 9110 747 9162 756
rect 9180 790 9232 799
rect 9180 756 9186 790
rect 9186 756 9220 790
rect 9220 756 9232 790
rect 9180 747 9232 756
rect 9250 790 9302 799
rect 9250 756 9259 790
rect 9259 756 9293 790
rect 9293 756 9302 790
rect 9250 747 9302 756
rect 9320 790 9372 799
rect 9320 756 9332 790
rect 9332 756 9366 790
rect 9366 756 9372 790
rect 9320 747 9372 756
rect 9558 790 9610 799
rect 9558 756 9564 790
rect 9564 756 9598 790
rect 9598 756 9610 790
rect 9558 747 9610 756
rect 9628 790 9680 799
rect 9628 756 9637 790
rect 9637 756 9671 790
rect 9671 756 9680 790
rect 9628 747 9680 756
rect 9698 790 9750 799
rect 9698 756 9710 790
rect 9710 756 9744 790
rect 9744 756 9750 790
rect 9698 747 9750 756
rect 9768 790 9820 799
rect 9768 756 9783 790
rect 9783 756 9817 790
rect 9817 756 9820 790
rect 9768 747 9820 756
rect 9838 790 9890 799
rect 9838 756 9856 790
rect 9856 756 9890 790
rect 9838 747 9890 756
rect 9908 790 9960 799
rect 9978 790 10030 799
rect 10048 790 10100 799
rect 10118 790 10170 799
rect 10189 790 10241 799
rect 10260 790 10312 799
rect 11558 797 11566 811
rect 11566 797 11600 811
rect 11600 797 11610 811
rect 9908 756 9929 790
rect 9929 756 9960 790
rect 9978 756 10002 790
rect 10002 756 10030 790
rect 10048 756 10075 790
rect 10075 756 10100 790
rect 10118 756 10148 790
rect 10148 756 10170 790
rect 10189 756 10221 790
rect 10221 756 10241 790
rect 10260 756 10294 790
rect 10294 756 10312 790
rect 9908 747 9960 756
rect 9978 747 10030 756
rect 10048 747 10100 756
rect 10118 747 10170 756
rect 10189 747 10241 756
rect 10260 747 10312 756
rect 11558 759 11610 797
rect 7322 723 7330 745
rect 7330 723 7364 745
rect 7364 723 7374 745
rect 7322 693 7374 723
rect 7322 649 7330 679
rect 7330 649 7364 679
rect 7364 649 7374 679
rect 7322 627 7374 649
rect 11558 723 11566 745
rect 11566 723 11600 745
rect 11600 723 11610 745
rect 11558 693 11610 723
rect 11558 649 11566 679
rect 11566 649 11600 679
rect 11600 649 11610 679
rect 7322 609 7374 613
rect 7322 575 7330 609
rect 7330 575 7364 609
rect 7364 575 7374 609
rect 7424 634 7476 643
rect 7496 634 7548 643
rect 7424 600 7454 634
rect 7454 600 7476 634
rect 7496 600 7528 634
rect 7528 600 7548 634
rect 7424 591 7476 600
rect 7496 591 7548 600
rect 7568 634 7620 643
rect 7568 600 7602 634
rect 7602 600 7620 634
rect 7568 591 7620 600
rect 7639 634 7691 643
rect 7639 600 7642 634
rect 7642 600 7676 634
rect 7676 600 7691 634
rect 7639 591 7691 600
rect 7710 634 7762 643
rect 7710 600 7716 634
rect 7716 600 7750 634
rect 7750 600 7762 634
rect 7710 591 7762 600
rect 7781 634 7833 643
rect 7781 600 7790 634
rect 7790 600 7824 634
rect 7824 600 7833 634
rect 7781 591 7833 600
rect 7852 634 7904 643
rect 7852 600 7864 634
rect 7864 600 7898 634
rect 7898 600 7904 634
rect 7852 591 7904 600
rect 7923 634 7975 643
rect 7923 600 7938 634
rect 7938 600 7972 634
rect 7972 600 7975 634
rect 7923 591 7975 600
rect 7994 634 8046 643
rect 7994 600 8012 634
rect 8012 600 8046 634
rect 7994 591 8046 600
rect 10458 634 10510 643
rect 10525 634 10577 643
rect 10591 634 10643 643
rect 10458 600 10474 634
rect 10474 600 10510 634
rect 10525 600 10548 634
rect 10548 600 10577 634
rect 10591 600 10622 634
rect 10622 600 10643 634
rect 10458 591 10510 600
rect 10525 591 10577 600
rect 10591 591 10643 600
rect 10657 634 10709 643
rect 10657 600 10662 634
rect 10662 600 10696 634
rect 10696 600 10709 634
rect 10657 591 10709 600
rect 10723 634 10775 643
rect 10723 600 10736 634
rect 10736 600 10770 634
rect 10770 600 10775 634
rect 10723 591 10775 600
rect 11558 627 11610 649
rect 11558 609 11610 613
rect 7322 561 7374 575
rect 7322 535 7374 547
rect 7322 501 7330 535
rect 7330 501 7364 535
rect 7364 501 7374 535
rect 7322 495 7374 501
rect 11558 575 11566 609
rect 11566 575 11600 609
rect 11600 575 11610 609
rect 11558 561 11610 575
rect 11558 535 11610 547
rect 11558 501 11566 535
rect 11566 501 11600 535
rect 11600 501 11610 535
rect 11558 495 11610 501
rect 8618 478 8670 487
rect 8689 478 8741 487
rect 8760 478 8812 487
rect 8830 478 8882 487
rect 8900 478 8952 487
rect 8970 478 9022 487
rect 8618 444 8636 478
rect 8636 444 8670 478
rect 8689 444 8709 478
rect 8709 444 8741 478
rect 8760 444 8782 478
rect 8782 444 8812 478
rect 8830 444 8855 478
rect 8855 444 8882 478
rect 8900 444 8928 478
rect 8928 444 8952 478
rect 8970 444 9001 478
rect 9001 444 9022 478
rect 8618 435 8670 444
rect 8689 435 8741 444
rect 8760 435 8812 444
rect 8830 435 8882 444
rect 8900 435 8952 444
rect 8970 435 9022 444
rect 9040 478 9092 487
rect 9040 444 9074 478
rect 9074 444 9092 478
rect 9040 435 9092 444
rect 9110 478 9162 487
rect 9110 444 9113 478
rect 9113 444 9147 478
rect 9147 444 9162 478
rect 9110 435 9162 444
rect 9180 478 9232 487
rect 9180 444 9186 478
rect 9186 444 9220 478
rect 9220 444 9232 478
rect 9180 435 9232 444
rect 9250 478 9302 487
rect 9250 444 9259 478
rect 9259 444 9293 478
rect 9293 444 9302 478
rect 9250 435 9302 444
rect 9320 478 9372 487
rect 9320 444 9332 478
rect 9332 444 9366 478
rect 9366 444 9372 478
rect 9320 435 9372 444
rect 9558 478 9610 487
rect 9558 444 9564 478
rect 9564 444 9598 478
rect 9598 444 9610 478
rect 9558 435 9610 444
rect 9628 478 9680 487
rect 9628 444 9637 478
rect 9637 444 9671 478
rect 9671 444 9680 478
rect 9628 435 9680 444
rect 9698 478 9750 487
rect 9698 444 9710 478
rect 9710 444 9744 478
rect 9744 444 9750 478
rect 9698 435 9750 444
rect 9768 478 9820 487
rect 9768 444 9783 478
rect 9783 444 9817 478
rect 9817 444 9820 478
rect 9768 435 9820 444
rect 9838 478 9890 487
rect 9838 444 9856 478
rect 9856 444 9890 478
rect 9838 435 9890 444
rect 9908 478 9960 487
rect 9978 478 10030 487
rect 10048 478 10100 487
rect 10118 478 10170 487
rect 10189 478 10241 487
rect 10260 478 10312 487
rect 9908 444 9929 478
rect 9929 444 9960 478
rect 9978 444 10002 478
rect 10002 444 10030 478
rect 10048 444 10075 478
rect 10075 444 10100 478
rect 10118 444 10148 478
rect 10148 444 10170 478
rect 10189 444 10221 478
rect 10221 444 10241 478
rect 10260 444 10294 478
rect 10294 444 10312 478
rect 9908 435 9960 444
rect 9978 435 10030 444
rect 10048 435 10100 444
rect 10118 435 10170 444
rect 10189 435 10241 444
rect 10260 435 10312 444
rect 8618 358 8670 383
rect 8684 358 8736 383
rect 8750 358 8802 383
rect 8816 358 8868 383
rect 8882 358 8934 383
rect 8948 358 9000 383
rect 9014 358 9066 383
rect 9080 358 9132 383
rect 9146 358 9198 383
rect 9212 358 9264 383
rect 9278 358 9330 383
rect 9344 358 9396 383
rect 9410 358 9462 383
rect 9476 358 9528 383
rect 9542 358 9594 383
rect 9608 358 9660 383
rect 9674 358 9726 383
rect 9740 358 9792 383
rect 9805 358 9857 383
rect 9870 358 9922 383
rect 9935 358 9987 383
rect 10000 358 10052 383
rect 10065 358 10117 383
rect 10130 358 10182 383
rect 10195 358 10247 383
rect 10260 358 10312 383
rect 8618 331 8670 358
rect 8684 331 8736 358
rect 8750 331 8802 358
rect 8816 331 8868 358
rect 8882 331 8934 358
rect 8948 331 9000 358
rect 9014 331 9066 358
rect 9080 331 9132 358
rect 9146 331 9198 358
rect 9212 331 9264 358
rect 9278 331 9330 358
rect 9344 331 9396 358
rect 9410 331 9462 358
rect 9476 331 9528 358
rect 9542 331 9594 358
rect 9608 331 9660 358
rect 9674 331 9726 358
rect 9740 331 9792 358
rect 9805 331 9857 358
rect 9870 331 9922 358
rect 9935 331 9987 358
rect 10000 331 10052 358
rect 10065 331 10117 358
rect 10130 331 10182 358
rect 10195 331 10247 358
rect 10260 331 10312 358
rect 7163 272 7215 324
rect 7229 286 7281 324
rect 7229 272 7235 286
rect 7235 272 7269 286
rect 7269 272 7281 286
rect 7295 286 7347 324
rect 7295 272 7308 286
rect 7308 272 7342 286
rect 7342 272 7347 286
rect 7361 286 7413 324
rect 7426 286 7478 324
rect 7491 286 7543 324
rect 7556 286 7608 324
rect 7621 286 7673 324
rect 7686 286 7738 324
rect 7751 286 7803 324
rect 7361 272 7381 286
rect 7381 272 7413 286
rect 7426 272 7454 286
rect 7454 272 7478 286
rect 7491 272 7527 286
rect 7527 272 7543 286
rect 7556 272 7561 286
rect 7561 272 7600 286
rect 7600 272 7608 286
rect 7621 272 7634 286
rect 7634 272 7673 286
rect 7686 272 7707 286
rect 7707 272 7738 286
rect 7751 272 7780 286
rect 7780 272 7803 286
rect 7816 286 7868 324
rect 7816 272 7819 286
rect 7819 272 7853 286
rect 7853 272 7868 286
rect 7881 286 7933 324
rect 7881 272 7892 286
rect 7892 272 7926 286
rect 7926 272 7933 286
rect 7946 286 7998 324
rect 8011 286 8063 324
rect 8076 286 8128 324
rect 7946 272 7965 286
rect 7965 272 7998 286
rect 8011 272 8038 286
rect 8038 272 8063 286
rect 8076 272 8111 286
rect 8111 272 8128 286
rect 7163 208 7215 260
rect 7229 252 7235 260
rect 7235 252 7269 260
rect 7269 252 7281 260
rect 7229 208 7281 252
rect 7295 252 7308 260
rect 7308 252 7342 260
rect 7342 252 7347 260
rect 7295 208 7347 252
rect 7361 252 7381 260
rect 7381 252 7413 260
rect 7426 252 7454 260
rect 7454 252 7478 260
rect 7491 252 7527 260
rect 7527 252 7543 260
rect 7556 252 7561 260
rect 7561 252 7600 260
rect 7600 252 7608 260
rect 7621 252 7634 260
rect 7634 252 7673 260
rect 7686 252 7707 260
rect 7707 252 7738 260
rect 7751 252 7780 260
rect 7780 252 7803 260
rect 7361 208 7413 252
rect 7426 208 7478 252
rect 7491 208 7543 252
rect 7556 208 7608 252
rect 7621 208 7673 252
rect 7686 208 7738 252
rect 7751 208 7803 252
rect 7816 252 7819 260
rect 7819 252 7853 260
rect 7853 252 7868 260
rect 7816 208 7868 252
rect 7881 252 7892 260
rect 7892 252 7926 260
rect 7926 252 7933 260
rect 7881 208 7933 252
rect 7946 252 7965 260
rect 7965 252 7998 260
rect 8011 252 8038 260
rect 8038 252 8063 260
rect 8076 252 8111 260
rect 8111 252 8128 260
rect 8618 267 8670 319
rect 8684 267 8736 319
rect 8750 267 8802 319
rect 8816 267 8868 319
rect 8882 267 8934 319
rect 8948 267 9000 319
rect 9014 267 9066 319
rect 9080 267 9132 319
rect 9146 267 9198 319
rect 9212 267 9264 319
rect 9278 267 9330 319
rect 9344 267 9396 319
rect 9410 267 9462 319
rect 9476 267 9528 319
rect 9542 267 9594 319
rect 9608 267 9660 319
rect 9674 267 9726 319
rect 9740 267 9792 319
rect 9805 267 9857 319
rect 9870 267 9922 319
rect 9935 267 9987 319
rect 10000 267 10052 319
rect 10065 267 10117 319
rect 10130 267 10182 319
rect 10195 267 10247 319
rect 10260 267 10312 319
rect 7946 208 7998 252
rect 8011 208 8063 252
rect 8076 208 8128 252
rect -195 -88 -150 -56
rect -150 -88 -143 -56
rect -131 -88 -116 -56
rect -116 -88 -79 -56
rect -195 -108 -143 -88
rect -131 -108 -79 -88
rect -195 -164 -143 -124
rect -131 -164 -79 -124
rect -195 -176 -150 -164
rect -150 -176 -143 -164
rect -131 -176 -116 -164
rect -116 -176 -79 -164
rect 5377 -281 5429 -229
rect 5441 -281 5493 -229
rect 5411 -1353 5463 -1301
rect 5411 -1417 5463 -1365
rect 5723 -1327 5775 -1301
rect 5846 -1270 5898 -1261
rect 5846 -1304 5852 -1270
rect 5852 -1304 5886 -1270
rect 5886 -1304 5898 -1270
rect 5846 -1313 5898 -1304
rect 5911 -1270 5963 -1261
rect 5911 -1304 5927 -1270
rect 5927 -1304 5961 -1270
rect 5961 -1304 5963 -1270
rect 5911 -1313 5963 -1304
rect 5976 -1270 6028 -1261
rect 6041 -1270 6093 -1261
rect 6106 -1270 6158 -1261
rect 6171 -1270 6223 -1261
rect 6236 -1270 6288 -1261
rect 5976 -1304 6002 -1270
rect 6002 -1304 6028 -1270
rect 6041 -1304 6077 -1270
rect 6077 -1304 6093 -1270
rect 6106 -1304 6111 -1270
rect 6111 -1304 6152 -1270
rect 6152 -1304 6158 -1270
rect 6171 -1304 6186 -1270
rect 6186 -1304 6223 -1270
rect 6236 -1304 6261 -1270
rect 6261 -1304 6288 -1270
rect 5976 -1313 6028 -1304
rect 6041 -1313 6093 -1304
rect 6106 -1313 6158 -1304
rect 6171 -1313 6223 -1304
rect 6236 -1313 6288 -1304
rect 6301 -1270 6353 -1261
rect 6301 -1304 6302 -1270
rect 6302 -1304 6336 -1270
rect 6336 -1304 6353 -1270
rect 6301 -1313 6353 -1304
rect 6365 -1270 6417 -1261
rect 6365 -1304 6377 -1270
rect 6377 -1304 6411 -1270
rect 6411 -1304 6417 -1270
rect 6365 -1313 6417 -1304
rect 6429 -1270 6481 -1261
rect 6493 -1270 6545 -1261
rect 6557 -1270 6609 -1261
rect 6621 -1270 6673 -1261
rect 6685 -1270 6737 -1261
rect 6429 -1304 6452 -1270
rect 6452 -1304 6481 -1270
rect 6493 -1304 6527 -1270
rect 6527 -1304 6545 -1270
rect 6557 -1304 6561 -1270
rect 6561 -1304 6602 -1270
rect 6602 -1304 6609 -1270
rect 6621 -1304 6636 -1270
rect 6636 -1304 6673 -1270
rect 6685 -1304 6710 -1270
rect 6710 -1304 6737 -1270
rect 6429 -1313 6481 -1304
rect 6493 -1313 6545 -1304
rect 6557 -1313 6609 -1304
rect 6621 -1313 6673 -1304
rect 6685 -1313 6737 -1304
rect 6749 -1270 6801 -1261
rect 6749 -1304 6750 -1270
rect 6750 -1304 6784 -1270
rect 6784 -1304 6801 -1270
rect 6749 -1313 6801 -1304
rect 6813 -1270 6865 -1261
rect 6813 -1304 6824 -1270
rect 6824 -1304 6858 -1270
rect 6858 -1304 6865 -1270
rect 6813 -1313 6865 -1304
rect 6877 -1270 6929 -1261
rect 6941 -1270 6993 -1261
rect 7005 -1270 7057 -1261
rect 7069 -1270 7121 -1261
rect 7133 -1270 7185 -1261
rect 7197 -1270 7249 -1261
rect 6877 -1304 6898 -1270
rect 6898 -1304 6929 -1270
rect 6941 -1304 6972 -1270
rect 6972 -1304 6993 -1270
rect 7005 -1304 7006 -1270
rect 7006 -1304 7046 -1270
rect 7046 -1304 7057 -1270
rect 7069 -1304 7080 -1270
rect 7080 -1304 7120 -1270
rect 7120 -1304 7121 -1270
rect 7133 -1304 7154 -1270
rect 7154 -1304 7185 -1270
rect 7197 -1304 7228 -1270
rect 7228 -1304 7249 -1270
rect 6877 -1313 6929 -1304
rect 6941 -1313 6993 -1304
rect 7005 -1313 7057 -1304
rect 7069 -1313 7121 -1304
rect 7133 -1313 7185 -1304
rect 7197 -1313 7249 -1304
rect 7261 -1270 7313 -1261
rect 7261 -1304 7268 -1270
rect 7268 -1304 7302 -1270
rect 7302 -1304 7313 -1270
rect 7261 -1313 7313 -1304
rect 7325 -1270 7377 -1261
rect 7325 -1304 7342 -1270
rect 7342 -1304 7376 -1270
rect 7376 -1304 7377 -1270
rect 7325 -1313 7377 -1304
rect 7389 -1270 7441 -1261
rect 7453 -1270 7505 -1261
rect 7517 -1270 7569 -1261
rect 7581 -1270 7633 -1261
rect 7645 -1270 7697 -1261
rect 7389 -1304 7416 -1270
rect 7416 -1304 7441 -1270
rect 7453 -1304 7490 -1270
rect 7490 -1304 7505 -1270
rect 7517 -1304 7524 -1270
rect 7524 -1304 7564 -1270
rect 7564 -1304 7569 -1270
rect 7581 -1304 7598 -1270
rect 7598 -1304 7633 -1270
rect 7645 -1304 7672 -1270
rect 7672 -1304 7697 -1270
rect 7389 -1313 7441 -1304
rect 7453 -1313 7505 -1304
rect 7517 -1313 7569 -1304
rect 7581 -1313 7633 -1304
rect 7645 -1313 7697 -1304
rect 7709 -1270 7761 -1261
rect 7709 -1304 7712 -1270
rect 7712 -1304 7746 -1270
rect 7746 -1304 7761 -1270
rect 7709 -1313 7761 -1304
rect 7773 -1270 7825 -1261
rect 7773 -1304 7786 -1270
rect 7786 -1304 7820 -1270
rect 7820 -1304 7825 -1270
rect 7773 -1313 7825 -1304
rect 5723 -1353 5734 -1327
rect 5734 -1353 5768 -1327
rect 5768 -1353 5775 -1327
rect 5723 -1399 5775 -1365
rect 5723 -1417 5734 -1399
rect 5734 -1417 5768 -1399
rect 5768 -1417 5775 -1399
rect 5846 -1426 5898 -1417
rect 5846 -1460 5852 -1426
rect 5852 -1460 5886 -1426
rect 5886 -1460 5898 -1426
rect 5846 -1469 5898 -1460
rect 5911 -1426 5963 -1417
rect 5911 -1460 5927 -1426
rect 5927 -1460 5961 -1426
rect 5961 -1460 5963 -1426
rect 5911 -1469 5963 -1460
rect 5976 -1426 6028 -1417
rect 6041 -1426 6093 -1417
rect 6106 -1426 6158 -1417
rect 6171 -1426 6223 -1417
rect 6236 -1426 6288 -1417
rect 5976 -1460 6002 -1426
rect 6002 -1460 6028 -1426
rect 6041 -1460 6077 -1426
rect 6077 -1460 6093 -1426
rect 6106 -1460 6111 -1426
rect 6111 -1460 6152 -1426
rect 6152 -1460 6158 -1426
rect 6171 -1460 6186 -1426
rect 6186 -1460 6223 -1426
rect 6236 -1460 6261 -1426
rect 6261 -1460 6288 -1426
rect 5976 -1469 6028 -1460
rect 6041 -1469 6093 -1460
rect 6106 -1469 6158 -1460
rect 6171 -1469 6223 -1460
rect 6236 -1469 6288 -1460
rect 6301 -1426 6353 -1417
rect 6301 -1460 6302 -1426
rect 6302 -1460 6336 -1426
rect 6336 -1460 6353 -1426
rect 6301 -1469 6353 -1460
rect 6365 -1426 6417 -1417
rect 6365 -1460 6377 -1426
rect 6377 -1460 6411 -1426
rect 6411 -1460 6417 -1426
rect 6365 -1469 6417 -1460
rect 6429 -1426 6481 -1417
rect 6493 -1426 6545 -1417
rect 6557 -1426 6609 -1417
rect 6621 -1426 6673 -1417
rect 6685 -1426 6737 -1417
rect 6429 -1460 6452 -1426
rect 6452 -1460 6481 -1426
rect 6493 -1460 6527 -1426
rect 6527 -1460 6545 -1426
rect 6557 -1460 6561 -1426
rect 6561 -1460 6602 -1426
rect 6602 -1460 6609 -1426
rect 6621 -1460 6636 -1426
rect 6636 -1460 6673 -1426
rect 6685 -1460 6710 -1426
rect 6710 -1460 6737 -1426
rect 6429 -1469 6481 -1460
rect 6493 -1469 6545 -1460
rect 6557 -1469 6609 -1460
rect 6621 -1469 6673 -1460
rect 6685 -1469 6737 -1460
rect 6749 -1426 6801 -1417
rect 6749 -1460 6750 -1426
rect 6750 -1460 6784 -1426
rect 6784 -1460 6801 -1426
rect 6749 -1469 6801 -1460
rect 6813 -1426 6865 -1417
rect 6813 -1460 6824 -1426
rect 6824 -1460 6858 -1426
rect 6858 -1460 6865 -1426
rect 6813 -1469 6865 -1460
rect 6877 -1426 6929 -1417
rect 6941 -1426 6993 -1417
rect 7005 -1426 7057 -1417
rect 7069 -1426 7121 -1417
rect 7133 -1426 7185 -1417
rect 7197 -1426 7249 -1417
rect 6877 -1460 6898 -1426
rect 6898 -1460 6929 -1426
rect 6941 -1460 6972 -1426
rect 6972 -1460 6993 -1426
rect 7005 -1460 7006 -1426
rect 7006 -1460 7046 -1426
rect 7046 -1460 7057 -1426
rect 7069 -1460 7080 -1426
rect 7080 -1460 7120 -1426
rect 7120 -1460 7121 -1426
rect 7133 -1460 7154 -1426
rect 7154 -1460 7185 -1426
rect 7197 -1460 7228 -1426
rect 7228 -1460 7249 -1426
rect 6877 -1469 6929 -1460
rect 6941 -1469 6993 -1460
rect 7005 -1469 7057 -1460
rect 7069 -1469 7121 -1460
rect 7133 -1469 7185 -1460
rect 7197 -1469 7249 -1460
rect 7261 -1426 7313 -1417
rect 7261 -1460 7268 -1426
rect 7268 -1460 7302 -1426
rect 7302 -1460 7313 -1426
rect 7261 -1469 7313 -1460
rect 7325 -1426 7377 -1417
rect 7325 -1460 7342 -1426
rect 7342 -1460 7376 -1426
rect 7376 -1460 7377 -1426
rect 7325 -1469 7377 -1460
rect 7389 -1426 7441 -1417
rect 7453 -1426 7505 -1417
rect 7517 -1426 7569 -1417
rect 7581 -1426 7633 -1417
rect 7645 -1426 7697 -1417
rect 7389 -1460 7416 -1426
rect 7416 -1460 7441 -1426
rect 7453 -1460 7490 -1426
rect 7490 -1460 7505 -1426
rect 7517 -1460 7524 -1426
rect 7524 -1460 7564 -1426
rect 7564 -1460 7569 -1426
rect 7581 -1460 7598 -1426
rect 7598 -1460 7633 -1426
rect 7645 -1460 7672 -1426
rect 7672 -1460 7697 -1426
rect 7389 -1469 7441 -1460
rect 7453 -1469 7505 -1460
rect 7517 -1469 7569 -1460
rect 7581 -1469 7633 -1460
rect 7645 -1469 7697 -1460
rect 7709 -1426 7761 -1417
rect 7709 -1460 7712 -1426
rect 7712 -1460 7746 -1426
rect 7746 -1460 7761 -1426
rect 7709 -1469 7761 -1460
rect 7773 -1426 7825 -1417
rect 7773 -1460 7786 -1426
rect 7786 -1460 7820 -1426
rect 7820 -1460 7825 -1426
rect 7773 -1469 7825 -1460
rect 5846 -1582 5898 -1573
rect 5846 -1616 5852 -1582
rect 5852 -1616 5886 -1582
rect 5886 -1616 5898 -1582
rect 5846 -1625 5898 -1616
rect 5911 -1582 5963 -1573
rect 5911 -1616 5927 -1582
rect 5927 -1616 5961 -1582
rect 5961 -1616 5963 -1582
rect 5911 -1625 5963 -1616
rect 5976 -1582 6028 -1573
rect 6041 -1582 6093 -1573
rect 6106 -1582 6158 -1573
rect 6171 -1582 6223 -1573
rect 6236 -1582 6288 -1573
rect 5976 -1616 6002 -1582
rect 6002 -1616 6028 -1582
rect 6041 -1616 6077 -1582
rect 6077 -1616 6093 -1582
rect 6106 -1616 6111 -1582
rect 6111 -1616 6152 -1582
rect 6152 -1616 6158 -1582
rect 6171 -1616 6186 -1582
rect 6186 -1616 6223 -1582
rect 6236 -1616 6261 -1582
rect 6261 -1616 6288 -1582
rect 5976 -1625 6028 -1616
rect 6041 -1625 6093 -1616
rect 6106 -1625 6158 -1616
rect 6171 -1625 6223 -1616
rect 6236 -1625 6288 -1616
rect 6301 -1582 6353 -1573
rect 6301 -1616 6302 -1582
rect 6302 -1616 6336 -1582
rect 6336 -1616 6353 -1582
rect 6301 -1625 6353 -1616
rect 6365 -1582 6417 -1573
rect 6365 -1616 6377 -1582
rect 6377 -1616 6411 -1582
rect 6411 -1616 6417 -1582
rect 6365 -1625 6417 -1616
rect 6429 -1582 6481 -1573
rect 6493 -1582 6545 -1573
rect 6557 -1582 6609 -1573
rect 6621 -1582 6673 -1573
rect 6685 -1582 6737 -1573
rect 6429 -1616 6452 -1582
rect 6452 -1616 6481 -1582
rect 6493 -1616 6527 -1582
rect 6527 -1616 6545 -1582
rect 6557 -1616 6561 -1582
rect 6561 -1616 6602 -1582
rect 6602 -1616 6609 -1582
rect 6621 -1616 6636 -1582
rect 6636 -1616 6673 -1582
rect 6685 -1616 6710 -1582
rect 6710 -1616 6737 -1582
rect 6429 -1625 6481 -1616
rect 6493 -1625 6545 -1616
rect 6557 -1625 6609 -1616
rect 6621 -1625 6673 -1616
rect 6685 -1625 6737 -1616
rect 6749 -1582 6801 -1573
rect 6749 -1616 6750 -1582
rect 6750 -1616 6784 -1582
rect 6784 -1616 6801 -1582
rect 6749 -1625 6801 -1616
rect 6813 -1582 6865 -1573
rect 6813 -1616 6824 -1582
rect 6824 -1616 6858 -1582
rect 6858 -1616 6865 -1582
rect 6813 -1625 6865 -1616
rect 6877 -1582 6929 -1573
rect 6941 -1582 6993 -1573
rect 7005 -1582 7057 -1573
rect 7069 -1582 7121 -1573
rect 7133 -1582 7185 -1573
rect 7197 -1582 7249 -1573
rect 6877 -1616 6898 -1582
rect 6898 -1616 6929 -1582
rect 6941 -1616 6972 -1582
rect 6972 -1616 6993 -1582
rect 7005 -1616 7006 -1582
rect 7006 -1616 7046 -1582
rect 7046 -1616 7057 -1582
rect 7069 -1616 7080 -1582
rect 7080 -1616 7120 -1582
rect 7120 -1616 7121 -1582
rect 7133 -1616 7154 -1582
rect 7154 -1616 7185 -1582
rect 7197 -1616 7228 -1582
rect 7228 -1616 7249 -1582
rect 6877 -1625 6929 -1616
rect 6941 -1625 6993 -1616
rect 7005 -1625 7057 -1616
rect 7069 -1625 7121 -1616
rect 7133 -1625 7185 -1616
rect 7197 -1625 7249 -1616
rect 7261 -1582 7313 -1573
rect 7261 -1616 7268 -1582
rect 7268 -1616 7302 -1582
rect 7302 -1616 7313 -1582
rect 7261 -1625 7313 -1616
rect 7325 -1582 7377 -1573
rect 7325 -1616 7342 -1582
rect 7342 -1616 7376 -1582
rect 7376 -1616 7377 -1582
rect 7325 -1625 7377 -1616
rect 7389 -1582 7441 -1573
rect 7453 -1582 7505 -1573
rect 7517 -1582 7569 -1573
rect 7581 -1582 7633 -1573
rect 7645 -1582 7697 -1573
rect 7389 -1616 7416 -1582
rect 7416 -1616 7441 -1582
rect 7453 -1616 7490 -1582
rect 7490 -1616 7505 -1582
rect 7517 -1616 7524 -1582
rect 7524 -1616 7564 -1582
rect 7564 -1616 7569 -1582
rect 7581 -1616 7598 -1582
rect 7598 -1616 7633 -1582
rect 7645 -1616 7672 -1582
rect 7672 -1616 7697 -1582
rect 7389 -1625 7441 -1616
rect 7453 -1625 7505 -1616
rect 7517 -1625 7569 -1616
rect 7581 -1625 7633 -1616
rect 7645 -1625 7697 -1616
rect 7709 -1582 7761 -1573
rect 7709 -1616 7712 -1582
rect 7712 -1616 7746 -1582
rect 7746 -1616 7761 -1582
rect 7709 -1625 7761 -1616
rect 7773 -1582 7825 -1573
rect 7773 -1616 7786 -1582
rect 7786 -1616 7820 -1582
rect 7820 -1616 7825 -1582
rect 7773 -1625 7825 -1616
rect 5846 -1738 5898 -1729
rect 5846 -1772 5852 -1738
rect 5852 -1772 5886 -1738
rect 5886 -1772 5898 -1738
rect 5846 -1781 5898 -1772
rect 5911 -1738 5963 -1729
rect 5911 -1772 5927 -1738
rect 5927 -1772 5961 -1738
rect 5961 -1772 5963 -1738
rect 5911 -1781 5963 -1772
rect 5976 -1738 6028 -1729
rect 6041 -1738 6093 -1729
rect 6106 -1738 6158 -1729
rect 6171 -1738 6223 -1729
rect 6236 -1738 6288 -1729
rect 5976 -1772 6002 -1738
rect 6002 -1772 6028 -1738
rect 6041 -1772 6077 -1738
rect 6077 -1772 6093 -1738
rect 6106 -1772 6111 -1738
rect 6111 -1772 6152 -1738
rect 6152 -1772 6158 -1738
rect 6171 -1772 6186 -1738
rect 6186 -1772 6223 -1738
rect 6236 -1772 6261 -1738
rect 6261 -1772 6288 -1738
rect 5976 -1781 6028 -1772
rect 6041 -1781 6093 -1772
rect 6106 -1781 6158 -1772
rect 6171 -1781 6223 -1772
rect 6236 -1781 6288 -1772
rect 6301 -1738 6353 -1729
rect 6301 -1772 6302 -1738
rect 6302 -1772 6336 -1738
rect 6336 -1772 6353 -1738
rect 6301 -1781 6353 -1772
rect 6365 -1738 6417 -1729
rect 6365 -1772 6377 -1738
rect 6377 -1772 6411 -1738
rect 6411 -1772 6417 -1738
rect 6365 -1781 6417 -1772
rect 6429 -1738 6481 -1729
rect 6493 -1738 6545 -1729
rect 6557 -1738 6609 -1729
rect 6621 -1738 6673 -1729
rect 6685 -1738 6737 -1729
rect 6429 -1772 6452 -1738
rect 6452 -1772 6481 -1738
rect 6493 -1772 6527 -1738
rect 6527 -1772 6545 -1738
rect 6557 -1772 6561 -1738
rect 6561 -1772 6602 -1738
rect 6602 -1772 6609 -1738
rect 6621 -1772 6636 -1738
rect 6636 -1772 6673 -1738
rect 6685 -1772 6710 -1738
rect 6710 -1772 6737 -1738
rect 6429 -1781 6481 -1772
rect 6493 -1781 6545 -1772
rect 6557 -1781 6609 -1772
rect 6621 -1781 6673 -1772
rect 6685 -1781 6737 -1772
rect 6749 -1738 6801 -1729
rect 6749 -1772 6750 -1738
rect 6750 -1772 6784 -1738
rect 6784 -1772 6801 -1738
rect 6749 -1781 6801 -1772
rect 6813 -1738 6865 -1729
rect 6813 -1772 6824 -1738
rect 6824 -1772 6858 -1738
rect 6858 -1772 6865 -1738
rect 6813 -1781 6865 -1772
rect 6877 -1738 6929 -1729
rect 6941 -1738 6993 -1729
rect 7005 -1738 7057 -1729
rect 7069 -1738 7121 -1729
rect 7133 -1738 7185 -1729
rect 7197 -1738 7249 -1729
rect 6877 -1772 6898 -1738
rect 6898 -1772 6929 -1738
rect 6941 -1772 6972 -1738
rect 6972 -1772 6993 -1738
rect 7005 -1772 7006 -1738
rect 7006 -1772 7046 -1738
rect 7046 -1772 7057 -1738
rect 7069 -1772 7080 -1738
rect 7080 -1772 7120 -1738
rect 7120 -1772 7121 -1738
rect 7133 -1772 7154 -1738
rect 7154 -1772 7185 -1738
rect 7197 -1772 7228 -1738
rect 7228 -1772 7249 -1738
rect 6877 -1781 6929 -1772
rect 6941 -1781 6993 -1772
rect 7005 -1781 7057 -1772
rect 7069 -1781 7121 -1772
rect 7133 -1781 7185 -1772
rect 7197 -1781 7249 -1772
rect 7261 -1738 7313 -1729
rect 7261 -1772 7268 -1738
rect 7268 -1772 7302 -1738
rect 7302 -1772 7313 -1738
rect 7261 -1781 7313 -1772
rect 7325 -1738 7377 -1729
rect 7325 -1772 7342 -1738
rect 7342 -1772 7376 -1738
rect 7376 -1772 7377 -1738
rect 7325 -1781 7377 -1772
rect 7389 -1738 7441 -1729
rect 7453 -1738 7505 -1729
rect 7517 -1738 7569 -1729
rect 7581 -1738 7633 -1729
rect 7645 -1738 7697 -1729
rect 7389 -1772 7416 -1738
rect 7416 -1772 7441 -1738
rect 7453 -1772 7490 -1738
rect 7490 -1772 7505 -1738
rect 7517 -1772 7524 -1738
rect 7524 -1772 7564 -1738
rect 7564 -1772 7569 -1738
rect 7581 -1772 7598 -1738
rect 7598 -1772 7633 -1738
rect 7645 -1772 7672 -1738
rect 7672 -1772 7697 -1738
rect 7389 -1781 7441 -1772
rect 7453 -1781 7505 -1772
rect 7517 -1781 7569 -1772
rect 7581 -1781 7633 -1772
rect 7645 -1781 7697 -1772
rect 7709 -1738 7761 -1729
rect 7709 -1772 7712 -1738
rect 7712 -1772 7746 -1738
rect 7746 -1772 7761 -1738
rect 7709 -1781 7761 -1772
rect 7773 -1738 7825 -1729
rect 7773 -1772 7786 -1738
rect 7786 -1772 7820 -1738
rect 7820 -1772 7825 -1738
rect 7773 -1781 7825 -1772
rect 7909 -1701 7961 -1692
rect 7909 -1735 7942 -1701
rect 7942 -1735 7961 -1701
rect 7909 -1744 7961 -1735
rect 7909 -1780 7961 -1766
rect 7909 -1814 7942 -1780
rect 7942 -1814 7961 -1780
rect 7909 -1818 7961 -1814
rect 5846 -1894 5898 -1885
rect 5846 -1928 5852 -1894
rect 5852 -1928 5886 -1894
rect 5886 -1928 5898 -1894
rect 5846 -1937 5898 -1928
rect 5911 -1894 5963 -1885
rect 5911 -1928 5927 -1894
rect 5927 -1928 5961 -1894
rect 5961 -1928 5963 -1894
rect 5911 -1937 5963 -1928
rect 5976 -1894 6028 -1885
rect 6041 -1894 6093 -1885
rect 6106 -1894 6158 -1885
rect 6171 -1894 6223 -1885
rect 6236 -1894 6288 -1885
rect 5976 -1928 6002 -1894
rect 6002 -1928 6028 -1894
rect 6041 -1928 6077 -1894
rect 6077 -1928 6093 -1894
rect 6106 -1928 6111 -1894
rect 6111 -1928 6152 -1894
rect 6152 -1928 6158 -1894
rect 6171 -1928 6186 -1894
rect 6186 -1928 6223 -1894
rect 6236 -1928 6261 -1894
rect 6261 -1928 6288 -1894
rect 5976 -1937 6028 -1928
rect 6041 -1937 6093 -1928
rect 6106 -1937 6158 -1928
rect 6171 -1937 6223 -1928
rect 6236 -1937 6288 -1928
rect 6301 -1894 6353 -1885
rect 6301 -1928 6302 -1894
rect 6302 -1928 6336 -1894
rect 6336 -1928 6353 -1894
rect 6301 -1937 6353 -1928
rect 6365 -1894 6417 -1885
rect 6365 -1928 6377 -1894
rect 6377 -1928 6411 -1894
rect 6411 -1928 6417 -1894
rect 6365 -1937 6417 -1928
rect 6429 -1894 6481 -1885
rect 6493 -1894 6545 -1885
rect 6557 -1894 6609 -1885
rect 6621 -1894 6673 -1885
rect 6685 -1894 6737 -1885
rect 6429 -1928 6452 -1894
rect 6452 -1928 6481 -1894
rect 6493 -1928 6527 -1894
rect 6527 -1928 6545 -1894
rect 6557 -1928 6561 -1894
rect 6561 -1928 6602 -1894
rect 6602 -1928 6609 -1894
rect 6621 -1928 6636 -1894
rect 6636 -1928 6673 -1894
rect 6685 -1928 6710 -1894
rect 6710 -1928 6737 -1894
rect 6429 -1937 6481 -1928
rect 6493 -1937 6545 -1928
rect 6557 -1937 6609 -1928
rect 6621 -1937 6673 -1928
rect 6685 -1937 6737 -1928
rect 6749 -1894 6801 -1885
rect 6749 -1928 6750 -1894
rect 6750 -1928 6784 -1894
rect 6784 -1928 6801 -1894
rect 6749 -1937 6801 -1928
rect 6813 -1894 6865 -1885
rect 6813 -1928 6824 -1894
rect 6824 -1928 6858 -1894
rect 6858 -1928 6865 -1894
rect 6813 -1937 6865 -1928
rect 6877 -1894 6929 -1885
rect 6941 -1894 6993 -1885
rect 7005 -1894 7057 -1885
rect 7069 -1894 7121 -1885
rect 7133 -1894 7185 -1885
rect 7197 -1894 7249 -1885
rect 6877 -1928 6898 -1894
rect 6898 -1928 6929 -1894
rect 6941 -1928 6972 -1894
rect 6972 -1928 6993 -1894
rect 7005 -1928 7006 -1894
rect 7006 -1928 7046 -1894
rect 7046 -1928 7057 -1894
rect 7069 -1928 7080 -1894
rect 7080 -1928 7120 -1894
rect 7120 -1928 7121 -1894
rect 7133 -1928 7154 -1894
rect 7154 -1928 7185 -1894
rect 7197 -1928 7228 -1894
rect 7228 -1928 7249 -1894
rect 6877 -1937 6929 -1928
rect 6941 -1937 6993 -1928
rect 7005 -1937 7057 -1928
rect 7069 -1937 7121 -1928
rect 7133 -1937 7185 -1928
rect 7197 -1937 7249 -1928
rect 7261 -1894 7313 -1885
rect 7261 -1928 7268 -1894
rect 7268 -1928 7302 -1894
rect 7302 -1928 7313 -1894
rect 7261 -1937 7313 -1928
rect 7325 -1894 7377 -1885
rect 7325 -1928 7342 -1894
rect 7342 -1928 7376 -1894
rect 7376 -1928 7377 -1894
rect 7325 -1937 7377 -1928
rect 7389 -1894 7441 -1885
rect 7453 -1894 7505 -1885
rect 7517 -1894 7569 -1885
rect 7581 -1894 7633 -1885
rect 7645 -1894 7697 -1885
rect 7389 -1928 7416 -1894
rect 7416 -1928 7441 -1894
rect 7453 -1928 7490 -1894
rect 7490 -1928 7505 -1894
rect 7517 -1928 7524 -1894
rect 7524 -1928 7564 -1894
rect 7564 -1928 7569 -1894
rect 7581 -1928 7598 -1894
rect 7598 -1928 7633 -1894
rect 7645 -1928 7672 -1894
rect 7672 -1928 7697 -1894
rect 7389 -1937 7441 -1928
rect 7453 -1937 7505 -1928
rect 7517 -1937 7569 -1928
rect 7581 -1937 7633 -1928
rect 7645 -1937 7697 -1928
rect 7709 -1894 7761 -1885
rect 7709 -1928 7712 -1894
rect 7712 -1928 7746 -1894
rect 7746 -1928 7761 -1894
rect 7709 -1937 7761 -1928
rect 7773 -1894 7825 -1885
rect 7773 -1928 7786 -1894
rect 7786 -1928 7820 -1894
rect 7820 -1928 7825 -1894
rect 7773 -1937 7825 -1928
rect 7909 -1859 7961 -1841
rect 7909 -1893 7942 -1859
rect 7942 -1893 7961 -1859
rect 7909 -1938 7961 -1916
rect 7909 -1968 7942 -1938
rect 7942 -1968 7961 -1938
rect 7909 -2043 7961 -1991
<< metal2 >>
rect -847 1736 11953 1856
rect -847 1582 -728 1736
tri -728 1701 -693 1736 nw
rect -679 1580 11953 1700
rect -679 1276 -558 1580
tri -558 1530 -508 1580 nw
tri 3103 1553 3130 1580 ne
rect -359 1494 -242 1500
rect -359 1442 -358 1494
rect -306 1442 -294 1494
rect -359 1421 -242 1442
rect -359 1369 -358 1421
rect -306 1369 -294 1421
rect -359 1348 -242 1369
rect -359 1296 -358 1348
rect -306 1296 -294 1348
rect -359 1267 -242 1296
tri -242 1267 -227 1282 sw
rect 3130 1267 3459 1580
tri 3459 1553 3486 1580 nw
rect -359 1215 -227 1267
tri -227 1215 -175 1267 sw
rect 3130 1215 3136 1267
rect 3188 1215 3203 1267
rect 3255 1215 3269 1267
rect 3321 1215 3335 1267
rect 3387 1215 3401 1267
rect 3453 1215 3459 1267
rect -359 1213 -175 1215
tri -175 1213 -173 1215 sw
rect -359 1212 -173 1213
tri -173 1212 -172 1213 sw
rect -359 1207 -172 1212
tri -172 1207 -167 1212 sw
rect 2305 1207 2361 1213
rect -359 1206 -167 1207
tri -167 1206 -166 1207 sw
tri -359 1155 -308 1206 ne
rect -308 1155 -166 1206
tri -166 1155 -115 1206 sw
rect 2357 1155 2361 1207
tri -308 1143 -296 1155 ne
rect -296 1143 -115 1155
tri -115 1143 -103 1155 sw
tri -296 1091 -244 1143 ne
rect -244 1091 640 1143
rect 692 1091 712 1143
rect 764 1091 784 1143
rect 836 1091 855 1143
rect 907 1091 913 1143
tri -244 1081 -234 1091 ne
rect -234 1081 913 1091
tri -234 1079 -232 1081 ne
rect -232 1079 913 1081
tri -232 1027 -180 1079 ne
rect -180 1027 640 1079
rect 692 1027 712 1079
rect 764 1027 784 1079
rect 836 1027 855 1079
rect 907 1027 913 1079
rect 1112 1141 2270 1147
rect 1112 1133 2154 1141
rect 1112 1081 1118 1133
rect 1170 1081 1195 1133
rect 1247 1081 1272 1133
rect 1324 1081 1348 1133
rect 1400 1081 1424 1133
rect 1476 1081 1500 1133
rect 1552 1089 2154 1133
rect 2206 1089 2218 1141
rect 1552 1081 2270 1089
rect 1112 1075 2270 1081
rect 1112 1055 2154 1075
rect 1112 1003 1118 1055
rect 1170 1003 1195 1055
rect 1247 1003 1272 1055
rect 1324 1003 1348 1055
rect 1400 1003 1424 1055
rect 1476 1003 1500 1055
rect 1552 1023 2154 1055
rect 2206 1023 2218 1075
rect 1552 1009 2270 1023
rect 1552 1003 2154 1009
rect 1112 997 2154 1003
tri 2108 973 2132 997 ne
rect 2132 973 2154 997
rect -509 967 436 973
rect -509 851 -490 967
rect -118 851 320 967
tri 2132 957 2148 973 ne
rect 2148 957 2154 973
rect 2206 957 2218 1009
tri 2148 951 2154 957 ne
rect 2154 951 2270 957
rect 2305 1134 2361 1155
rect 2357 1082 2361 1134
rect 2305 1061 2361 1082
rect 2357 1009 2361 1061
rect 2305 988 2361 1009
rect -509 845 436 851
rect 2357 936 2361 988
rect 2305 915 2361 936
rect 2357 863 2361 915
rect 2305 842 2361 863
tri -47 744 5 796 se
rect 5 744 640 796
rect 692 744 712 796
rect 764 744 784 796
rect 836 744 855 796
rect 907 744 913 796
tri -59 732 -47 744 se
rect -47 732 913 744
tri -79 712 -59 732 se
rect -59 712 640 732
rect -79 680 640 712
rect 692 680 712 732
rect 764 680 784 732
rect 836 680 855 732
rect 907 680 913 732
rect 2357 790 2361 842
rect 2305 769 2361 790
rect 2357 717 2361 769
rect 3130 955 3459 1215
rect 3130 903 3136 955
rect 3188 903 3203 955
rect 3255 903 3269 955
rect 3321 903 3335 955
rect 3387 903 3401 955
rect 3453 903 3459 955
rect 3130 756 3459 903
rect 3593 1404 3599 1456
rect 3651 1404 3665 1456
rect 3717 1404 3731 1456
rect 3783 1404 3797 1456
rect 3849 1404 3863 1456
rect 3915 1404 3929 1456
rect 3981 1404 3995 1456
rect 4047 1404 4061 1456
rect 4113 1404 4127 1456
rect 4179 1404 4193 1456
rect 4245 1404 4259 1456
rect 4311 1404 4325 1456
rect 4377 1404 4391 1456
rect 4443 1404 4457 1456
rect 4509 1404 4523 1456
rect 4575 1404 4589 1456
rect 4641 1404 4655 1456
rect 4707 1404 4721 1456
rect 4773 1404 4786 1456
rect 4838 1404 4851 1456
rect 4903 1404 4916 1456
rect 4968 1404 4981 1456
rect 5033 1404 5046 1456
rect 5098 1404 5111 1456
rect 5163 1404 5176 1456
rect 5228 1404 5241 1456
rect 5293 1404 5299 1456
rect 3593 1392 5299 1404
rect 3593 1340 3599 1392
rect 3651 1340 3665 1392
rect 3717 1340 3731 1392
rect 3783 1340 3797 1392
rect 3849 1340 3863 1392
rect 3915 1340 3929 1392
rect 3981 1340 3995 1392
rect 4047 1340 4061 1392
rect 4113 1340 4127 1392
rect 4179 1340 4193 1392
rect 4245 1340 4259 1392
rect 4311 1340 4325 1392
rect 4377 1340 4391 1392
rect 4443 1340 4457 1392
rect 4509 1340 4523 1392
rect 4575 1340 4589 1392
rect 4641 1340 4655 1392
rect 4707 1340 4721 1392
rect 4773 1340 4786 1392
rect 4838 1340 4851 1392
rect 4903 1340 4916 1392
rect 4968 1340 4981 1392
rect 5033 1340 5046 1392
rect 5098 1340 5111 1392
rect 5163 1340 5176 1392
rect 5228 1340 5241 1392
rect 5293 1340 5299 1392
rect 3593 1111 5299 1340
rect 6644 1450 6895 1456
rect 6696 1447 6716 1450
rect 6768 1447 6788 1450
rect 6840 1447 6895 1450
rect 6644 1391 6679 1398
rect 6735 1391 6759 1398
rect 6815 1391 6839 1398
rect 6644 1379 6895 1391
rect 6696 1365 6716 1379
rect 6768 1365 6788 1379
rect 6840 1365 6895 1379
rect 6644 1309 6679 1327
rect 6735 1309 6759 1327
rect 6815 1309 6839 1327
rect 6644 1300 6895 1309
rect 8612 1404 8618 1456
rect 8670 1404 8684 1456
rect 8736 1404 8750 1456
rect 8802 1404 8816 1456
rect 8868 1404 8882 1456
rect 8934 1404 8948 1456
rect 9000 1404 9014 1456
rect 9066 1404 9080 1456
rect 9132 1404 9146 1456
rect 9198 1404 9212 1456
rect 9264 1404 9278 1456
rect 9330 1404 9344 1456
rect 9396 1404 9410 1456
rect 9462 1404 9476 1456
rect 9528 1404 9542 1456
rect 9594 1404 9608 1456
rect 9660 1404 9674 1456
rect 9726 1404 9740 1456
rect 9792 1404 9805 1456
rect 9857 1404 9870 1456
rect 9922 1404 9935 1456
rect 9987 1404 10000 1456
rect 10052 1404 10065 1456
rect 10117 1404 10130 1456
rect 10182 1404 10195 1456
rect 10247 1404 10260 1456
rect 10312 1404 10318 1456
rect 8612 1392 10318 1404
rect 8612 1340 8618 1392
rect 8670 1340 8684 1392
rect 8736 1340 8750 1392
rect 8802 1340 8816 1392
rect 8868 1340 8882 1392
rect 8934 1340 8948 1392
rect 9000 1340 9014 1392
rect 9066 1340 9080 1392
rect 9132 1340 9146 1392
rect 9198 1340 9212 1392
rect 9264 1340 9278 1392
rect 9330 1340 9344 1392
rect 9396 1340 9410 1392
rect 9462 1340 9476 1392
rect 9528 1340 9542 1392
rect 9594 1340 9608 1392
rect 9660 1340 9674 1392
rect 9726 1340 9740 1392
rect 9792 1340 9805 1392
rect 9857 1340 9870 1392
rect 9922 1340 9935 1392
rect 9987 1340 10000 1392
rect 10052 1340 10065 1392
rect 10117 1340 10130 1392
rect 10182 1340 10195 1392
rect 10247 1340 10260 1392
rect 10312 1340 10318 1392
rect 5814 1267 5823 1269
rect 5879 1267 5904 1269
rect 5960 1267 5984 1269
rect 6040 1267 6064 1269
rect 6120 1267 6144 1269
rect 6200 1267 6224 1269
rect 6280 1267 6304 1269
rect 6360 1267 6384 1269
rect 6440 1267 6455 1269
rect 5814 1215 5820 1267
rect 5879 1215 5885 1267
rect 6129 1215 6141 1267
rect 6200 1215 6205 1267
rect 6449 1215 6455 1267
rect 5814 1213 5823 1215
rect 5879 1213 5904 1215
rect 5960 1213 5984 1215
rect 6040 1213 6064 1215
rect 6120 1213 6144 1215
rect 6200 1213 6224 1215
rect 6280 1213 6304 1215
rect 6360 1213 6384 1215
rect 6440 1213 6455 1215
rect 6539 1264 7374 1272
rect 6591 1212 7374 1264
rect 7418 1267 7427 1269
rect 7483 1267 7507 1269
rect 7563 1267 7587 1269
rect 7643 1267 7667 1269
rect 7723 1267 7747 1269
rect 7803 1267 7827 1269
rect 7883 1267 7907 1269
rect 7963 1267 7987 1269
rect 8043 1267 8052 1269
rect 7418 1215 7424 1267
rect 7483 1215 7496 1267
rect 7563 1215 7568 1267
rect 7904 1215 7907 1267
rect 7975 1215 7987 1267
rect 8046 1215 8052 1267
rect 7418 1213 7427 1215
rect 7483 1213 7507 1215
rect 7563 1213 7587 1215
rect 7643 1213 7667 1215
rect 7723 1213 7747 1215
rect 7803 1213 7827 1215
rect 7883 1213 7907 1215
rect 7963 1213 7987 1215
rect 8043 1213 8052 1215
rect 6539 1207 7374 1212
rect 6539 1195 7322 1207
rect 6539 1191 6613 1195
rect 6591 1155 6613 1191
tri 6613 1155 6653 1195 nw
tri 7259 1155 7299 1195 ne
rect 7299 1155 7322 1195
rect 6591 1141 6599 1155
tri 6599 1141 6613 1155 nw
tri 7299 1141 7313 1155 ne
rect 7313 1141 7374 1155
rect 6539 1133 6591 1139
tri 6591 1133 6599 1141 nw
tri 7313 1136 7318 1141 ne
tri 6672 1111 6674 1113 se
rect 6674 1111 6683 1113
rect 3593 1059 3599 1111
rect 3651 1059 3670 1111
rect 3722 1059 3741 1111
rect 3793 1059 3811 1111
rect 3863 1059 3881 1111
rect 3933 1059 3951 1111
rect 4003 1059 4021 1111
rect 4073 1059 4091 1111
rect 4143 1059 4161 1111
rect 4213 1059 4231 1111
rect 4283 1059 4301 1111
rect 4353 1059 4539 1111
rect 4591 1059 4609 1111
rect 4661 1059 4679 1111
rect 4731 1059 4749 1111
rect 4801 1059 4819 1111
rect 4871 1059 4889 1111
rect 4941 1059 4959 1111
rect 5011 1059 5029 1111
rect 5081 1059 5099 1111
rect 5151 1059 5170 1111
rect 5222 1059 5241 1111
rect 5293 1059 5299 1111
rect 3593 799 5299 1059
rect 6156 1059 6162 1111
rect 6214 1059 6250 1111
rect 6302 1059 6338 1111
rect 6390 1100 6399 1111
tri 6399 1100 6410 1111 sw
tri 6661 1100 6672 1111 se
rect 6672 1100 6683 1111
rect 6390 1059 6683 1100
rect 6156 1057 6683 1059
rect 6739 1057 6766 1113
rect 6822 1057 6849 1113
rect 6905 1057 6914 1113
rect 7318 1089 7322 1141
rect 7318 1075 7374 1089
rect 6156 1044 6698 1057
tri 6698 1044 6711 1057 nw
rect 7318 1023 7322 1075
rect 7318 1009 7374 1023
rect 7318 957 7322 1009
rect 8612 1111 10318 1340
rect 10452 1267 10461 1269
rect 10517 1267 10546 1269
rect 10602 1267 10631 1269
rect 10687 1267 10716 1269
rect 10772 1267 10781 1269
rect 10452 1215 10458 1267
rect 10517 1215 10525 1267
rect 10709 1215 10716 1267
rect 10775 1215 10781 1267
rect 10452 1213 10461 1215
rect 10517 1213 10546 1215
rect 10602 1213 10631 1215
rect 10687 1213 10716 1215
rect 10772 1213 10781 1215
rect 8612 1059 8618 1111
rect 8670 1059 8689 1111
rect 8741 1059 8760 1111
rect 8812 1059 8830 1111
rect 8882 1059 8900 1111
rect 8952 1059 8970 1111
rect 9022 1059 9040 1111
rect 9092 1059 9110 1111
rect 9162 1059 9180 1111
rect 9232 1059 9250 1111
rect 9302 1059 9320 1111
rect 9372 1059 9558 1111
rect 9610 1059 9628 1111
rect 9680 1059 9698 1111
rect 9750 1059 9768 1111
rect 9820 1059 9838 1111
rect 9890 1059 9908 1111
rect 9960 1059 9978 1111
rect 10030 1059 10048 1111
rect 10100 1059 10118 1111
rect 10170 1059 10189 1111
rect 10241 1059 10260 1111
rect 10312 1059 10318 1111
rect 5814 955 5823 957
rect 5879 955 5904 957
rect 5960 955 5984 957
rect 6040 955 6064 957
rect 6120 955 6144 957
rect 6200 955 6224 957
rect 6280 955 6304 957
rect 6360 955 6384 957
rect 6440 955 6455 957
rect 5814 903 5820 955
rect 5879 903 5885 955
rect 6129 903 6141 955
rect 6200 903 6205 955
rect 6449 903 6455 955
rect 5814 901 5823 903
rect 5879 901 5904 903
rect 5960 901 5984 903
rect 6040 901 6064 903
rect 6120 901 6144 903
rect 6200 901 6224 903
rect 6280 901 6304 903
rect 6360 901 6384 903
rect 6440 901 6455 903
rect 7318 943 7374 957
rect 7318 891 7322 943
rect 7418 955 7427 957
rect 7483 955 7520 957
rect 7576 955 7612 957
rect 7668 955 7704 957
rect 7760 955 7796 957
rect 7852 955 7888 957
rect 7944 955 7980 957
rect 8036 955 8045 957
rect 7418 903 7424 955
rect 7483 903 7495 955
rect 7689 903 7704 955
rect 7760 903 7777 955
rect 7969 903 7980 955
rect 8039 903 8045 955
rect 7418 901 7427 903
rect 7483 901 7520 903
rect 7576 901 7612 903
rect 7668 901 7704 903
rect 7760 901 7796 903
rect 7852 901 7888 903
rect 7944 901 7980 903
rect 8036 901 8045 903
rect 7318 877 7374 891
rect 7318 825 7322 877
rect 7318 811 7374 825
tri 6672 799 6674 801 se
rect 6674 799 6683 801
rect 2305 697 2361 717
tri -195 -50 -79 66 se
rect -79 -50 37 680
tri 37 645 72 680 nw
rect 1111 630 1117 682
rect 1169 630 1194 682
rect 1246 630 1271 682
rect 1323 630 1348 682
rect 1400 630 1424 682
rect 1476 630 1500 682
rect 1552 630 1558 682
rect 1111 604 1558 630
rect 467 598 519 604
rect 467 534 519 546
rect 467 212 519 482
rect 1111 552 1117 604
rect 1169 552 1194 604
rect 1246 552 1271 604
rect 1323 552 1348 604
rect 1400 552 1424 604
rect 1476 552 1500 604
rect 1552 552 1558 604
rect 1111 362 1558 552
rect 2357 645 2361 697
rect 3593 747 3599 799
rect 3651 747 3670 799
rect 3722 747 3741 799
rect 3793 747 3811 799
rect 3863 747 3881 799
rect 3933 747 3951 799
rect 4003 747 4021 799
rect 4073 747 4091 799
rect 4143 747 4161 799
rect 4213 747 4231 799
rect 4283 747 4301 799
rect 4353 747 4539 799
rect 4591 747 4609 799
rect 4661 747 4679 799
rect 4731 747 4749 799
rect 4801 747 4819 799
rect 4871 747 4889 799
rect 4941 747 4959 799
rect 5011 747 5029 799
rect 5081 747 5099 799
rect 5151 747 5170 799
rect 5222 747 5241 799
rect 5293 747 5299 799
rect 6156 747 6162 799
rect 6214 747 6250 799
rect 6302 747 6338 799
rect 6390 747 6683 799
tri 1558 362 1573 377 sw
rect 1111 340 1573 362
tri 1573 340 1595 362 sw
rect 1111 331 1595 340
tri 1595 331 1604 340 sw
rect 1111 324 1604 331
tri 1604 324 1611 331 sw
rect 1111 276 1611 324
tri 1611 276 1659 324 sw
rect 2305 323 2361 645
rect 3130 643 3459 688
rect 3130 591 3136 643
rect 3188 591 3203 643
rect 3255 591 3269 643
rect 3321 591 3335 643
rect 3387 591 3401 643
rect 3453 591 3459 643
rect 3130 438 3459 591
rect 3593 487 5299 747
tri 6672 745 6674 747 ne
rect 6674 745 6683 747
rect 6739 745 6766 801
rect 6822 745 6849 801
rect 6905 745 6914 801
rect 7318 759 7322 811
rect 7318 745 7374 759
rect 6535 704 6591 710
tri 6526 657 6535 666 se
rect 6535 657 6539 704
rect 6526 652 6539 657
rect 7318 693 7322 745
rect 7318 679 7374 693
tri 6591 657 6600 666 sw
rect 6591 652 6600 657
rect 5814 643 5823 645
rect 5879 643 5904 645
rect 5960 643 5984 645
rect 6040 643 6064 645
rect 6120 643 6144 645
rect 6200 643 6224 645
rect 6280 643 6304 645
rect 6360 643 6384 645
rect 6440 643 6455 645
rect 5814 591 5820 643
rect 5879 591 5885 643
rect 6129 591 6141 643
rect 6200 591 6205 643
rect 6449 591 6455 643
rect 5814 589 5823 591
rect 5879 589 5904 591
rect 5960 589 5984 591
rect 6040 589 6064 591
rect 6120 589 6144 591
rect 6200 589 6224 591
rect 6280 589 6304 591
rect 6360 589 6384 591
rect 6440 589 6455 591
rect 6526 634 6600 652
rect 6526 578 6535 634
rect 6591 578 6600 634
rect 6526 554 6600 578
rect 6526 498 6535 554
rect 6591 498 6600 554
rect 6526 489 6600 498
rect 7318 627 7322 679
rect 8612 799 10318 1059
rect 11554 1207 11610 1213
rect 11554 1155 11558 1207
rect 11554 1141 11610 1155
rect 11554 1089 11558 1141
rect 11554 1075 11610 1089
rect 11554 1023 11558 1075
rect 11554 1009 11610 1023
rect 11554 957 11558 1009
rect 10452 955 10461 957
rect 10517 955 10546 957
rect 10602 955 10631 957
rect 10687 955 10716 957
rect 10772 955 10781 957
rect 10452 903 10458 955
rect 10517 903 10525 955
rect 10709 903 10716 955
rect 10775 903 10781 955
rect 10452 901 10461 903
rect 10517 901 10546 903
rect 10602 901 10631 903
rect 10687 901 10716 903
rect 10772 901 10781 903
rect 11554 943 11610 957
rect 8612 747 8618 799
rect 8670 747 8689 799
rect 8741 747 8760 799
rect 8812 747 8830 799
rect 8882 747 8900 799
rect 8952 747 8970 799
rect 9022 747 9040 799
rect 9092 747 9110 799
rect 9162 747 9180 799
rect 9232 747 9250 799
rect 9302 747 9320 799
rect 9372 747 9558 799
rect 9610 747 9628 799
rect 9680 747 9698 799
rect 9750 747 9768 799
rect 9820 747 9838 799
rect 9890 747 9908 799
rect 9960 747 9978 799
rect 10030 747 10048 799
rect 10100 747 10118 799
rect 10170 747 10189 799
rect 10241 747 10260 799
rect 10312 747 10318 799
rect 7318 613 7374 627
rect 7318 561 7322 613
rect 7418 643 7427 645
rect 7483 643 7507 645
rect 7563 643 7587 645
rect 7643 643 7667 645
rect 7723 643 7747 645
rect 7803 643 7827 645
rect 7883 643 7907 645
rect 7963 643 7987 645
rect 8043 643 8052 645
rect 7418 591 7424 643
rect 7483 591 7496 643
rect 7563 591 7568 643
rect 7904 591 7907 643
rect 7975 591 7987 643
rect 8046 591 8052 643
rect 7418 589 7427 591
rect 7483 589 7507 591
rect 7563 589 7587 591
rect 7643 589 7667 591
rect 7723 589 7747 591
rect 7803 589 7827 591
rect 7883 589 7907 591
rect 7963 589 7987 591
rect 8043 589 8052 591
rect 7318 547 7374 561
rect 7318 495 7322 547
rect 7318 489 7374 495
rect 3593 435 3599 487
rect 3651 435 3670 487
rect 3722 435 3741 487
rect 3793 435 3811 487
rect 3863 435 3881 487
rect 3933 435 3951 487
rect 4003 435 4021 487
rect 4073 435 4091 487
rect 4143 435 4161 487
rect 4213 435 4231 487
rect 4283 435 4301 487
rect 4353 435 4539 487
rect 4591 435 4609 487
rect 4661 435 4679 487
rect 4731 435 4749 487
rect 4801 435 4819 487
rect 4871 435 4889 487
rect 4941 435 4959 487
rect 5011 435 5029 487
rect 5081 435 5099 487
rect 5151 435 5170 487
rect 5222 435 5241 487
rect 5293 435 5299 487
rect 8612 487 10318 747
rect 11554 891 11558 943
rect 11554 877 11610 891
rect 11554 825 11558 877
rect 11554 811 11610 825
rect 11554 759 11558 811
rect 11554 745 11610 759
rect 11554 693 11558 745
rect 11554 679 11610 693
rect 10452 643 10461 645
rect 10517 643 10546 645
rect 10602 643 10631 645
rect 10687 643 10716 645
rect 10772 643 10781 645
rect 10452 591 10458 643
rect 10517 591 10525 643
rect 10709 591 10716 643
rect 10775 591 10781 643
rect 10452 589 10461 591
rect 10517 589 10546 591
rect 10602 589 10631 591
rect 10687 589 10716 591
rect 10772 589 10781 591
rect 11554 627 11558 679
rect 11554 613 11610 627
tri 6664 456 6687 479 se
rect 6687 470 6903 479
rect 3593 414 5299 435
rect 3593 362 3599 414
rect 3651 362 3665 414
rect 3717 362 3731 414
rect 3783 362 3797 414
rect 3849 362 3863 414
rect 3915 362 3929 414
rect 3981 362 3995 414
rect 4047 362 4061 414
rect 4113 362 4127 414
rect 4179 362 4193 414
rect 4245 362 4259 414
rect 4311 362 4325 414
rect 4377 362 4391 414
rect 4443 362 4457 414
rect 4509 362 4523 414
rect 4575 362 4589 414
rect 4641 362 4655 414
rect 4707 362 4721 414
rect 4773 362 4786 414
rect 4838 362 4851 414
rect 4903 362 4916 414
rect 4968 362 4981 414
rect 5033 362 5046 414
rect 5098 362 5111 414
rect 5163 362 5176 414
rect 5228 362 5241 414
rect 5293 362 5299 414
rect 6177 340 6183 456
rect 6363 414 6687 456
rect 6743 414 6767 470
rect 6823 414 6847 470
rect 6363 388 6903 414
rect 6363 340 6687 388
tri 6670 331 6679 340 ne
rect 6679 332 6687 340
rect 6743 332 6767 388
rect 6823 332 6847 388
rect 8612 435 8618 487
rect 8670 435 8689 487
rect 8741 435 8760 487
rect 8812 435 8830 487
rect 8882 435 8900 487
rect 8952 435 8970 487
rect 9022 435 9040 487
rect 9092 435 9110 487
rect 9162 435 9180 487
rect 9232 435 9250 487
rect 9302 435 9320 487
rect 9372 435 9558 487
rect 9610 435 9628 487
rect 9680 435 9698 487
rect 9750 435 9768 487
rect 9820 435 9838 487
rect 9890 435 9908 487
rect 9960 435 9978 487
rect 10030 435 10048 487
rect 10100 435 10118 487
rect 10170 435 10189 487
rect 10241 435 10260 487
rect 10312 435 10318 487
tri 7106 383 7107 384 se
rect 7107 383 8383 384
tri 8383 383 8384 384 sw
rect 8612 383 10318 435
tri 7096 373 7106 383 se
rect 7106 373 8384 383
tri 8384 373 8394 383 sw
rect 6679 331 6903 332
tri 7054 331 7096 373 se
rect 7096 352 8394 373
rect 7096 331 7114 352
tri 7114 331 7135 352 nw
tri 8334 331 8355 352 ne
rect 8355 331 8394 352
tri 8394 331 8436 373 sw
rect 8612 331 8618 383
rect 8670 331 8684 383
rect 8736 331 8750 383
rect 8802 331 8816 383
rect 8868 331 8882 383
rect 8934 331 8948 383
rect 9000 331 9014 383
rect 9066 331 9080 383
rect 9132 331 9146 383
rect 9198 331 9212 383
rect 9264 331 9278 383
rect 9330 331 9344 383
rect 9396 331 9410 383
rect 9462 331 9476 383
rect 9528 331 9542 383
rect 9594 331 9608 383
rect 9660 331 9674 383
rect 9726 331 9740 383
rect 9792 331 9805 383
rect 9857 331 9870 383
rect 9922 331 9935 383
rect 9987 331 10000 383
rect 10052 331 10065 383
rect 10117 331 10130 383
rect 10182 331 10195 383
rect 10247 331 10260 383
rect 10312 331 10318 383
tri 6679 324 6686 331 ne
rect 6686 324 6903 331
tri 7047 324 7054 331 se
rect 7054 324 7107 331
tri 7107 324 7114 331 nw
tri 8355 324 8362 331 ne
rect 8362 324 8436 331
tri 2361 323 2362 324 sw
tri 6686 323 6687 324 ne
rect 6687 323 6903 324
tri 7046 323 7047 324 se
rect 7047 323 7075 324
rect 2305 304 2362 323
tri 2362 304 2381 323 sw
tri 7027 304 7046 323 se
rect 7046 304 7075 323
rect 2305 288 2381 304
tri 2381 288 2397 304 sw
tri 4749 288 4765 304 se
rect 4765 292 4932 304
tri 4932 292 4944 304 sw
tri 7015 292 7027 304 se
rect 7027 292 7075 304
tri 7075 292 7107 324 nw
rect 4765 288 4944 292
rect 2305 280 3494 288
tri 3494 280 3502 288 sw
tri 4741 280 4749 288 se
rect 4749 280 4944 288
tri 4944 280 4956 292 sw
tri 7003 280 7015 292 se
rect 7015 280 7063 292
tri 7063 280 7075 292 nw
rect 2305 276 7059 280
tri 7059 276 7063 280 nw
rect 1111 272 1659 276
tri 1659 272 1663 276 sw
rect 2305 272 7055 276
tri 7055 272 7059 276 nw
rect 7157 272 7163 324
rect 7215 272 7229 324
rect 7281 272 7295 324
rect 7347 272 7361 324
rect 7413 272 7426 324
rect 7478 272 7491 324
rect 7543 272 7556 324
rect 7608 272 7621 324
rect 7673 272 7686 324
rect 7738 272 7751 324
rect 7803 272 7816 324
rect 7868 272 7881 324
rect 7933 272 7946 324
rect 7998 272 8011 324
rect 8063 272 8076 324
rect 8128 272 8134 324
tri 8362 319 8367 324 ne
rect 8367 323 8436 324
tri 8436 323 8444 331 sw
rect 8367 319 8444 323
tri 8444 319 8448 323 sw
rect 8612 319 10318 331
tri 8367 292 8394 319 ne
rect 8394 292 8448 319
tri 8448 292 8475 319 sw
tri 8394 280 8406 292 ne
rect 8406 280 8475 292
tri 8406 276 8410 280 ne
rect 8410 276 8475 280
tri 8475 276 8491 292 sw
rect 1111 267 1663 272
tri 1663 267 1668 272 sw
rect 2305 267 7050 272
tri 7050 267 7055 272 nw
rect 1111 260 1668 267
tri 1668 260 1675 267 sw
rect 2305 260 7043 267
tri 7043 260 7050 267 nw
rect 7157 260 8134 272
tri 8410 267 8419 276 ne
rect 8419 267 8491 276
tri 8491 267 8500 276 sw
rect 8612 267 8618 319
rect 8670 267 8684 319
rect 8736 267 8750 319
rect 8802 267 8816 319
rect 8868 267 8882 319
rect 8934 267 8948 319
rect 9000 267 9014 319
rect 9066 267 9080 319
rect 9132 267 9146 319
rect 9198 267 9212 319
rect 9264 267 9278 319
rect 9330 267 9344 319
rect 9396 267 9410 319
rect 9462 267 9476 319
rect 9528 267 9542 319
rect 9594 267 9608 319
rect 9660 267 9674 319
rect 9726 267 9740 319
rect 9792 267 9805 319
rect 9857 267 9870 319
rect 9922 267 9935 319
rect 9987 267 10000 319
rect 10052 267 10065 319
rect 10117 267 10130 319
rect 10182 267 10195 319
rect 10247 267 10260 319
rect 10312 267 10318 319
rect 11554 561 11558 613
rect 11554 547 11610 561
rect 11554 495 11558 547
tri 11545 267 11554 276 se
rect 11554 267 11610 495
rect 1111 256 1675 260
tri 1675 256 1679 260 sw
rect 2305 256 7039 260
tri 7039 256 7043 260 nw
rect 1111 228 1679 256
tri 1679 228 1707 256 sw
tri 3467 248 3475 256 ne
rect 3475 248 7031 256
tri 7031 248 7039 256 nw
tri 7149 248 7157 256 se
rect 7157 248 7163 260
tri 7129 228 7149 248 se
rect 7149 228 7163 248
rect 1111 220 1707 228
tri 1707 220 1715 228 sw
tri 7121 220 7129 228 se
rect 7129 220 7163 228
rect 1111 208 7163 220
rect 7215 208 7229 260
rect 7281 208 7295 260
rect 7347 208 7361 260
rect 7413 208 7426 260
rect 7478 208 7491 260
rect 7543 208 7556 260
rect 7608 208 7621 260
rect 7673 208 7686 260
rect 7738 208 7751 260
rect 7803 208 7816 260
rect 7868 208 7881 260
rect 7933 208 7946 260
rect 7998 208 8011 260
rect 8063 208 8076 260
rect 8128 208 8134 260
tri 8419 256 8430 267 ne
rect 8430 256 8500 267
tri 8500 256 8511 267 sw
tri 11534 256 11545 267 se
rect 11545 256 11610 267
tri 8430 220 8466 256 ne
rect 8466 228 8511 256
tri 8511 228 8539 256 sw
tri 11506 228 11534 256 se
rect 11534 228 11610 256
rect 8466 220 8539 228
tri 8539 220 8547 228 sw
tri 10399 220 10407 228 se
rect 10407 220 11610 228
tri 8466 211 8475 220 ne
rect 8475 211 8547 220
tri 8547 211 8556 220 sw
tri 10390 211 10399 220 se
rect 10399 211 11610 220
rect 1111 140 8134 208
tri 8475 201 8485 211 ne
rect 8485 201 11610 211
tri 8485 179 8507 201 ne
rect 8507 196 11610 201
rect 8507 179 10439 196
tri 10439 179 10456 196 nw
rect -195 -56 37 -50
rect -143 -108 -131 -56
rect -79 -108 37 -56
rect -195 -124 37 -108
rect -143 -176 -131 -124
rect -79 -176 37 -124
rect -195 -182 37 -176
rect 5371 -281 5377 -229
rect 5429 -281 5441 -229
rect 5493 -281 5499 -229
rect 5411 -1301 5775 -1293
rect 5463 -1353 5723 -1301
rect 5820 -1315 5829 -1259
rect 5885 -1261 5921 -1259
rect 5977 -1261 6013 -1259
rect 6069 -1261 6105 -1259
rect 6161 -1261 6197 -1259
rect 6253 -1261 6289 -1259
rect 6345 -1261 6380 -1259
rect 6436 -1261 6445 -1259
rect 7238 -1261 7247 -1259
rect 7303 -1261 7335 -1259
rect 7391 -1261 7422 -1259
rect 7478 -1261 7509 -1259
rect 7565 -1261 7596 -1259
rect 7652 -1261 7683 -1259
rect 7739 -1261 7770 -1259
rect 5898 -1313 5911 -1261
rect 6093 -1313 6105 -1261
rect 6161 -1313 6171 -1261
rect 6288 -1313 6289 -1261
rect 6353 -1313 6365 -1261
rect 6481 -1313 6493 -1261
rect 6545 -1313 6557 -1261
rect 6609 -1313 6621 -1261
rect 6673 -1313 6685 -1261
rect 6737 -1313 6749 -1261
rect 6801 -1313 6813 -1261
rect 6865 -1313 6877 -1261
rect 6929 -1313 6941 -1261
rect 6993 -1313 7005 -1261
rect 7057 -1313 7069 -1261
rect 7121 -1313 7133 -1261
rect 7185 -1313 7197 -1261
rect 7313 -1313 7325 -1261
rect 7505 -1313 7509 -1261
rect 7569 -1313 7581 -1261
rect 7761 -1313 7770 -1261
rect 5885 -1315 5921 -1313
rect 5977 -1315 6013 -1313
rect 6069 -1315 6105 -1313
rect 6161 -1315 6197 -1313
rect 6253 -1315 6289 -1313
rect 6345 -1315 6380 -1313
rect 6436 -1315 6445 -1313
rect 7238 -1315 7247 -1313
rect 7303 -1315 7335 -1313
rect 7391 -1315 7422 -1313
rect 7478 -1315 7509 -1313
rect 7565 -1315 7596 -1313
rect 7652 -1315 7683 -1313
rect 7739 -1315 7770 -1313
rect 7826 -1315 7835 -1259
rect 5411 -1365 5775 -1353
rect 5463 -1417 5723 -1365
rect 6670 -1417 6679 -1415
rect 6735 -1417 6766 -1415
rect 6822 -1417 6853 -1415
rect 6909 -1417 6918 -1415
rect 5411 -1423 5775 -1417
rect 5840 -1469 5846 -1417
rect 5898 -1469 5911 -1417
rect 5963 -1469 5976 -1417
rect 6028 -1469 6041 -1417
rect 6093 -1469 6106 -1417
rect 6158 -1469 6171 -1417
rect 6223 -1469 6236 -1417
rect 6288 -1469 6301 -1417
rect 6353 -1469 6365 -1417
rect 6417 -1469 6429 -1417
rect 6481 -1469 6493 -1417
rect 6545 -1469 6557 -1417
rect 6609 -1469 6621 -1417
rect 6673 -1469 6679 -1417
rect 6737 -1469 6749 -1417
rect 6929 -1469 6941 -1417
rect 6993 -1469 7005 -1417
rect 7057 -1469 7069 -1417
rect 7121 -1469 7133 -1417
rect 7185 -1469 7197 -1417
rect 7249 -1469 7261 -1417
rect 7313 -1469 7325 -1417
rect 7377 -1469 7389 -1417
rect 7441 -1469 7453 -1417
rect 7505 -1469 7517 -1417
rect 7569 -1469 7581 -1417
rect 7633 -1469 7645 -1417
rect 7697 -1469 7709 -1417
rect 7761 -1469 7773 -1417
rect 7825 -1469 7831 -1417
rect 6670 -1471 6679 -1469
rect 6735 -1471 6766 -1469
rect 6822 -1471 6853 -1469
rect 6909 -1471 6918 -1469
rect 5820 -1627 5829 -1571
rect 5885 -1573 5921 -1571
rect 5977 -1573 6013 -1571
rect 6069 -1573 6105 -1571
rect 6161 -1573 6197 -1571
rect 6253 -1573 6289 -1571
rect 6345 -1573 6380 -1571
rect 6436 -1573 6445 -1571
rect 7238 -1573 7247 -1571
rect 7303 -1573 7335 -1571
rect 7391 -1573 7422 -1571
rect 7478 -1573 7509 -1571
rect 7565 -1573 7596 -1571
rect 7652 -1573 7683 -1571
rect 7739 -1573 7770 -1571
rect 5898 -1625 5911 -1573
rect 6093 -1625 6105 -1573
rect 6161 -1625 6171 -1573
rect 6288 -1625 6289 -1573
rect 6353 -1625 6365 -1573
rect 6481 -1625 6493 -1573
rect 6545 -1625 6557 -1573
rect 6609 -1625 6621 -1573
rect 6673 -1625 6685 -1573
rect 6737 -1625 6749 -1573
rect 6801 -1625 6813 -1573
rect 6865 -1625 6877 -1573
rect 6929 -1625 6941 -1573
rect 6993 -1625 7005 -1573
rect 7057 -1625 7069 -1573
rect 7121 -1625 7133 -1573
rect 7185 -1625 7197 -1573
rect 7313 -1625 7325 -1573
rect 7505 -1625 7509 -1573
rect 7569 -1625 7581 -1573
rect 7761 -1625 7770 -1573
rect 5885 -1627 5921 -1625
rect 5977 -1627 6013 -1625
rect 6069 -1627 6105 -1625
rect 6161 -1627 6197 -1625
rect 6253 -1627 6289 -1625
rect 6345 -1627 6380 -1625
rect 6436 -1627 6445 -1625
rect 7238 -1627 7247 -1625
rect 7303 -1627 7335 -1625
rect 7391 -1627 7422 -1625
rect 7478 -1627 7509 -1625
rect 7565 -1627 7596 -1625
rect 7652 -1627 7683 -1625
rect 7739 -1627 7770 -1625
rect 7826 -1627 7835 -1571
rect 7890 -1692 7980 -1686
rect 6670 -1729 6679 -1727
rect 6735 -1729 6766 -1727
rect 6822 -1729 6853 -1727
rect 6909 -1729 6918 -1727
rect 5840 -1781 5846 -1729
rect 5898 -1781 5911 -1729
rect 5963 -1781 5976 -1729
rect 6028 -1781 6041 -1729
rect 6093 -1781 6106 -1729
rect 6158 -1781 6171 -1729
rect 6223 -1781 6236 -1729
rect 6288 -1781 6301 -1729
rect 6353 -1781 6365 -1729
rect 6417 -1781 6429 -1729
rect 6481 -1781 6493 -1729
rect 6545 -1781 6557 -1729
rect 6609 -1781 6621 -1729
rect 6673 -1781 6679 -1729
rect 6737 -1781 6749 -1729
rect 6929 -1781 6941 -1729
rect 6993 -1781 7005 -1729
rect 7057 -1781 7069 -1729
rect 7121 -1781 7133 -1729
rect 7185 -1781 7197 -1729
rect 7249 -1781 7261 -1729
rect 7313 -1781 7325 -1729
rect 7377 -1781 7389 -1729
rect 7441 -1781 7453 -1729
rect 7505 -1781 7517 -1729
rect 7569 -1781 7581 -1729
rect 7633 -1781 7645 -1729
rect 7697 -1781 7709 -1729
rect 7761 -1781 7773 -1729
rect 7825 -1781 7831 -1729
rect 7890 -1744 7909 -1692
rect 7961 -1744 7980 -1692
rect 7890 -1766 7980 -1744
rect 6670 -1783 6679 -1781
rect 6735 -1783 6766 -1781
rect 6822 -1783 6853 -1781
rect 6909 -1783 6918 -1781
rect 7890 -1818 7909 -1766
rect 7961 -1818 7980 -1766
rect 7890 -1841 7980 -1818
rect 5820 -1939 5829 -1883
rect 5885 -1885 5921 -1883
rect 5977 -1885 6013 -1883
rect 6069 -1885 6105 -1883
rect 6161 -1885 6197 -1883
rect 6253 -1885 6289 -1883
rect 6345 -1885 6380 -1883
rect 6436 -1885 6445 -1883
rect 7238 -1885 7247 -1883
rect 7303 -1885 7335 -1883
rect 7391 -1885 7422 -1883
rect 7478 -1885 7509 -1883
rect 7565 -1885 7596 -1883
rect 7652 -1885 7683 -1883
rect 7739 -1885 7770 -1883
rect 5898 -1937 5911 -1885
rect 6093 -1937 6105 -1885
rect 6161 -1937 6171 -1885
rect 6288 -1937 6289 -1885
rect 6353 -1937 6365 -1885
rect 6481 -1937 6493 -1885
rect 6545 -1937 6557 -1885
rect 6609 -1937 6621 -1885
rect 6673 -1937 6685 -1885
rect 6737 -1937 6749 -1885
rect 6801 -1937 6813 -1885
rect 6865 -1937 6877 -1885
rect 6929 -1937 6941 -1885
rect 6993 -1937 7005 -1885
rect 7057 -1937 7069 -1885
rect 7121 -1937 7133 -1885
rect 7185 -1937 7197 -1885
rect 7313 -1937 7325 -1885
rect 7505 -1937 7509 -1885
rect 7569 -1937 7581 -1885
rect 7761 -1937 7770 -1885
rect 5885 -1939 5921 -1937
rect 5977 -1939 6013 -1937
rect 6069 -1939 6105 -1937
rect 6161 -1939 6197 -1937
rect 6253 -1939 6289 -1937
rect 6345 -1939 6380 -1937
rect 6436 -1939 6445 -1937
rect 7238 -1939 7247 -1937
rect 7303 -1939 7335 -1937
rect 7391 -1939 7422 -1937
rect 7478 -1939 7509 -1937
rect 7565 -1939 7596 -1937
rect 7652 -1939 7683 -1937
rect 7739 -1939 7770 -1937
rect 7826 -1939 7835 -1883
rect 7890 -1893 7909 -1841
rect 7961 -1893 7980 -1841
rect 7890 -1916 7980 -1893
rect 7890 -1968 7909 -1916
rect 7961 -1968 7980 -1916
rect 7890 -1991 7980 -1968
rect 7890 -2043 7909 -1991
rect 7961 -2043 7980 -1991
rect 7890 -2049 7980 -2043
rect 6535 -2686 6605 -2677
rect 6591 -2742 6605 -2686
rect 6535 -2766 6605 -2742
rect 6591 -2822 6605 -2766
rect 6535 -2831 6605 -2822
<< via2 >>
rect 6679 1398 6696 1447
rect 6696 1398 6716 1447
rect 6716 1398 6735 1447
rect 6759 1398 6768 1447
rect 6768 1398 6788 1447
rect 6788 1398 6815 1447
rect 6839 1398 6840 1447
rect 6840 1398 6895 1447
rect 6679 1391 6735 1398
rect 6759 1391 6815 1398
rect 6839 1391 6895 1398
rect 6679 1327 6696 1365
rect 6696 1327 6716 1365
rect 6716 1327 6735 1365
rect 6759 1327 6768 1365
rect 6768 1327 6788 1365
rect 6788 1327 6815 1365
rect 6839 1327 6840 1365
rect 6840 1327 6895 1365
rect 6679 1309 6735 1327
rect 6759 1309 6815 1327
rect 6839 1309 6895 1327
rect 5823 1267 5879 1269
rect 5904 1267 5960 1269
rect 5984 1267 6040 1269
rect 6064 1267 6120 1269
rect 6144 1267 6200 1269
rect 6224 1267 6280 1269
rect 6304 1267 6360 1269
rect 6384 1267 6440 1269
rect 5823 1215 5872 1267
rect 5872 1215 5879 1267
rect 5904 1215 5937 1267
rect 5937 1215 5949 1267
rect 5949 1215 5960 1267
rect 5984 1215 6001 1267
rect 6001 1215 6013 1267
rect 6013 1215 6040 1267
rect 6064 1215 6065 1267
rect 6065 1215 6077 1267
rect 6077 1215 6120 1267
rect 6144 1215 6193 1267
rect 6193 1215 6200 1267
rect 6224 1215 6257 1267
rect 6257 1215 6269 1267
rect 6269 1215 6280 1267
rect 6304 1215 6321 1267
rect 6321 1215 6333 1267
rect 6333 1215 6360 1267
rect 6384 1215 6385 1267
rect 6385 1215 6397 1267
rect 6397 1215 6440 1267
rect 5823 1213 5879 1215
rect 5904 1213 5960 1215
rect 5984 1213 6040 1215
rect 6064 1213 6120 1215
rect 6144 1213 6200 1215
rect 6224 1213 6280 1215
rect 6304 1213 6360 1215
rect 6384 1213 6440 1215
rect 7427 1267 7483 1269
rect 7507 1267 7563 1269
rect 7587 1267 7643 1269
rect 7667 1267 7723 1269
rect 7747 1267 7803 1269
rect 7827 1267 7883 1269
rect 7907 1267 7963 1269
rect 7987 1267 8043 1269
rect 7427 1215 7476 1267
rect 7476 1215 7483 1267
rect 7507 1215 7548 1267
rect 7548 1215 7563 1267
rect 7587 1215 7620 1267
rect 7620 1215 7639 1267
rect 7639 1215 7643 1267
rect 7667 1215 7691 1267
rect 7691 1215 7710 1267
rect 7710 1215 7723 1267
rect 7747 1215 7762 1267
rect 7762 1215 7781 1267
rect 7781 1215 7803 1267
rect 7827 1215 7833 1267
rect 7833 1215 7852 1267
rect 7852 1215 7883 1267
rect 7907 1215 7923 1267
rect 7923 1215 7963 1267
rect 7987 1215 7994 1267
rect 7994 1215 8043 1267
rect 7427 1213 7483 1215
rect 7507 1213 7563 1215
rect 7587 1213 7643 1215
rect 7667 1213 7723 1215
rect 7747 1213 7803 1215
rect 7827 1213 7883 1215
rect 7907 1213 7963 1215
rect 7987 1213 8043 1215
rect 6683 1057 6739 1113
rect 6766 1057 6822 1113
rect 6849 1057 6905 1113
rect 10461 1267 10517 1269
rect 10546 1267 10602 1269
rect 10631 1267 10687 1269
rect 10716 1267 10772 1269
rect 10461 1215 10510 1267
rect 10510 1215 10517 1267
rect 10546 1215 10577 1267
rect 10577 1215 10591 1267
rect 10591 1215 10602 1267
rect 10631 1215 10643 1267
rect 10643 1215 10657 1267
rect 10657 1215 10687 1267
rect 10716 1215 10723 1267
rect 10723 1215 10772 1267
rect 10461 1213 10517 1215
rect 10546 1213 10602 1215
rect 10631 1213 10687 1215
rect 10716 1213 10772 1215
rect 5823 955 5879 957
rect 5904 955 5960 957
rect 5984 955 6040 957
rect 6064 955 6120 957
rect 6144 955 6200 957
rect 6224 955 6280 957
rect 6304 955 6360 957
rect 6384 955 6440 957
rect 5823 903 5872 955
rect 5872 903 5879 955
rect 5904 903 5937 955
rect 5937 903 5949 955
rect 5949 903 5960 955
rect 5984 903 6001 955
rect 6001 903 6013 955
rect 6013 903 6040 955
rect 6064 903 6065 955
rect 6065 903 6077 955
rect 6077 903 6120 955
rect 6144 903 6193 955
rect 6193 903 6200 955
rect 6224 903 6257 955
rect 6257 903 6269 955
rect 6269 903 6280 955
rect 6304 903 6321 955
rect 6321 903 6333 955
rect 6333 903 6360 955
rect 6384 903 6385 955
rect 6385 903 6397 955
rect 6397 903 6440 955
rect 5823 901 5879 903
rect 5904 901 5960 903
rect 5984 901 6040 903
rect 6064 901 6120 903
rect 6144 901 6200 903
rect 6224 901 6280 903
rect 6304 901 6360 903
rect 6384 901 6440 903
rect 7427 955 7483 957
rect 7520 955 7576 957
rect 7612 955 7668 957
rect 7704 955 7760 957
rect 7796 955 7852 957
rect 7888 955 7944 957
rect 7980 955 8036 957
rect 7427 903 7476 955
rect 7476 903 7483 955
rect 7520 903 7547 955
rect 7547 903 7566 955
rect 7566 903 7576 955
rect 7612 903 7618 955
rect 7618 903 7637 955
rect 7637 903 7668 955
rect 7704 903 7707 955
rect 7707 903 7759 955
rect 7759 903 7760 955
rect 7796 903 7829 955
rect 7829 903 7847 955
rect 7847 903 7852 955
rect 7888 903 7899 955
rect 7899 903 7917 955
rect 7917 903 7944 955
rect 7980 903 7987 955
rect 7987 903 8036 955
rect 7427 901 7483 903
rect 7520 901 7576 903
rect 7612 901 7668 903
rect 7704 901 7760 903
rect 7796 901 7852 903
rect 7888 901 7944 903
rect 7980 901 8036 903
rect 6683 745 6739 801
rect 6766 745 6822 801
rect 6849 745 6905 801
rect 5823 643 5879 645
rect 5904 643 5960 645
rect 5984 643 6040 645
rect 6064 643 6120 645
rect 6144 643 6200 645
rect 6224 643 6280 645
rect 6304 643 6360 645
rect 6384 643 6440 645
rect 5823 591 5872 643
rect 5872 591 5879 643
rect 5904 591 5937 643
rect 5937 591 5949 643
rect 5949 591 5960 643
rect 5984 591 6001 643
rect 6001 591 6013 643
rect 6013 591 6040 643
rect 6064 591 6065 643
rect 6065 591 6077 643
rect 6077 591 6120 643
rect 6144 591 6193 643
rect 6193 591 6200 643
rect 6224 591 6257 643
rect 6257 591 6269 643
rect 6269 591 6280 643
rect 6304 591 6321 643
rect 6321 591 6333 643
rect 6333 591 6360 643
rect 6384 591 6385 643
rect 6385 591 6397 643
rect 6397 591 6440 643
rect 5823 589 5879 591
rect 5904 589 5960 591
rect 5984 589 6040 591
rect 6064 589 6120 591
rect 6144 589 6200 591
rect 6224 589 6280 591
rect 6304 589 6360 591
rect 6384 589 6440 591
rect 6535 631 6591 634
rect 6535 579 6539 631
rect 6539 579 6591 631
rect 6535 578 6591 579
rect 6535 498 6591 554
rect 10461 955 10517 957
rect 10546 955 10602 957
rect 10631 955 10687 957
rect 10716 955 10772 957
rect 10461 903 10510 955
rect 10510 903 10517 955
rect 10546 903 10577 955
rect 10577 903 10591 955
rect 10591 903 10602 955
rect 10631 903 10643 955
rect 10643 903 10657 955
rect 10657 903 10687 955
rect 10716 903 10723 955
rect 10723 903 10772 955
rect 10461 901 10517 903
rect 10546 901 10602 903
rect 10631 901 10687 903
rect 10716 901 10772 903
rect 7427 643 7483 645
rect 7507 643 7563 645
rect 7587 643 7643 645
rect 7667 643 7723 645
rect 7747 643 7803 645
rect 7827 643 7883 645
rect 7907 643 7963 645
rect 7987 643 8043 645
rect 7427 591 7476 643
rect 7476 591 7483 643
rect 7507 591 7548 643
rect 7548 591 7563 643
rect 7587 591 7620 643
rect 7620 591 7639 643
rect 7639 591 7643 643
rect 7667 591 7691 643
rect 7691 591 7710 643
rect 7710 591 7723 643
rect 7747 591 7762 643
rect 7762 591 7781 643
rect 7781 591 7803 643
rect 7827 591 7833 643
rect 7833 591 7852 643
rect 7852 591 7883 643
rect 7907 591 7923 643
rect 7923 591 7963 643
rect 7987 591 7994 643
rect 7994 591 8043 643
rect 7427 589 7483 591
rect 7507 589 7563 591
rect 7587 589 7643 591
rect 7667 589 7723 591
rect 7747 589 7803 591
rect 7827 589 7883 591
rect 7907 589 7963 591
rect 7987 589 8043 591
rect 10461 643 10517 645
rect 10546 643 10602 645
rect 10631 643 10687 645
rect 10716 643 10772 645
rect 10461 591 10510 643
rect 10510 591 10517 643
rect 10546 591 10577 643
rect 10577 591 10591 643
rect 10591 591 10602 643
rect 10631 591 10643 643
rect 10643 591 10657 643
rect 10657 591 10687 643
rect 10716 591 10723 643
rect 10723 591 10772 643
rect 10461 589 10517 591
rect 10546 589 10602 591
rect 10631 589 10687 591
rect 10716 589 10772 591
rect 6687 414 6743 470
rect 6767 414 6823 470
rect 6847 414 6903 470
rect 6687 332 6743 388
rect 6767 332 6823 388
rect 6847 332 6903 388
rect 5829 -1261 5885 -1259
rect 5921 -1261 5977 -1259
rect 6013 -1261 6069 -1259
rect 6105 -1261 6161 -1259
rect 6197 -1261 6253 -1259
rect 6289 -1261 6345 -1259
rect 6380 -1261 6436 -1259
rect 7247 -1261 7303 -1259
rect 7335 -1261 7391 -1259
rect 7422 -1261 7478 -1259
rect 7509 -1261 7565 -1259
rect 7596 -1261 7652 -1259
rect 7683 -1261 7739 -1259
rect 7770 -1261 7826 -1259
rect 5829 -1313 5846 -1261
rect 5846 -1313 5885 -1261
rect 5921 -1313 5963 -1261
rect 5963 -1313 5976 -1261
rect 5976 -1313 5977 -1261
rect 6013 -1313 6028 -1261
rect 6028 -1313 6041 -1261
rect 6041 -1313 6069 -1261
rect 6105 -1313 6106 -1261
rect 6106 -1313 6158 -1261
rect 6158 -1313 6161 -1261
rect 6197 -1313 6223 -1261
rect 6223 -1313 6236 -1261
rect 6236 -1313 6253 -1261
rect 6289 -1313 6301 -1261
rect 6301 -1313 6345 -1261
rect 6380 -1313 6417 -1261
rect 6417 -1313 6429 -1261
rect 6429 -1313 6436 -1261
rect 7247 -1313 7249 -1261
rect 7249 -1313 7261 -1261
rect 7261 -1313 7303 -1261
rect 7335 -1313 7377 -1261
rect 7377 -1313 7389 -1261
rect 7389 -1313 7391 -1261
rect 7422 -1313 7441 -1261
rect 7441 -1313 7453 -1261
rect 7453 -1313 7478 -1261
rect 7509 -1313 7517 -1261
rect 7517 -1313 7565 -1261
rect 7596 -1313 7633 -1261
rect 7633 -1313 7645 -1261
rect 7645 -1313 7652 -1261
rect 7683 -1313 7697 -1261
rect 7697 -1313 7709 -1261
rect 7709 -1313 7739 -1261
rect 7770 -1313 7773 -1261
rect 7773 -1313 7825 -1261
rect 7825 -1313 7826 -1261
rect 5829 -1315 5885 -1313
rect 5921 -1315 5977 -1313
rect 6013 -1315 6069 -1313
rect 6105 -1315 6161 -1313
rect 6197 -1315 6253 -1313
rect 6289 -1315 6345 -1313
rect 6380 -1315 6436 -1313
rect 7247 -1315 7303 -1313
rect 7335 -1315 7391 -1313
rect 7422 -1315 7478 -1313
rect 7509 -1315 7565 -1313
rect 7596 -1315 7652 -1313
rect 7683 -1315 7739 -1313
rect 7770 -1315 7826 -1313
rect 6679 -1417 6735 -1415
rect 6766 -1417 6822 -1415
rect 6853 -1417 6909 -1415
rect 6679 -1469 6685 -1417
rect 6685 -1469 6735 -1417
rect 6766 -1469 6801 -1417
rect 6801 -1469 6813 -1417
rect 6813 -1469 6822 -1417
rect 6853 -1469 6865 -1417
rect 6865 -1469 6877 -1417
rect 6877 -1469 6909 -1417
rect 6679 -1471 6735 -1469
rect 6766 -1471 6822 -1469
rect 6853 -1471 6909 -1469
rect 5829 -1573 5885 -1571
rect 5921 -1573 5977 -1571
rect 6013 -1573 6069 -1571
rect 6105 -1573 6161 -1571
rect 6197 -1573 6253 -1571
rect 6289 -1573 6345 -1571
rect 6380 -1573 6436 -1571
rect 7247 -1573 7303 -1571
rect 7335 -1573 7391 -1571
rect 7422 -1573 7478 -1571
rect 7509 -1573 7565 -1571
rect 7596 -1573 7652 -1571
rect 7683 -1573 7739 -1571
rect 7770 -1573 7826 -1571
rect 5829 -1625 5846 -1573
rect 5846 -1625 5885 -1573
rect 5921 -1625 5963 -1573
rect 5963 -1625 5976 -1573
rect 5976 -1625 5977 -1573
rect 6013 -1625 6028 -1573
rect 6028 -1625 6041 -1573
rect 6041 -1625 6069 -1573
rect 6105 -1625 6106 -1573
rect 6106 -1625 6158 -1573
rect 6158 -1625 6161 -1573
rect 6197 -1625 6223 -1573
rect 6223 -1625 6236 -1573
rect 6236 -1625 6253 -1573
rect 6289 -1625 6301 -1573
rect 6301 -1625 6345 -1573
rect 6380 -1625 6417 -1573
rect 6417 -1625 6429 -1573
rect 6429 -1625 6436 -1573
rect 7247 -1625 7249 -1573
rect 7249 -1625 7261 -1573
rect 7261 -1625 7303 -1573
rect 7335 -1625 7377 -1573
rect 7377 -1625 7389 -1573
rect 7389 -1625 7391 -1573
rect 7422 -1625 7441 -1573
rect 7441 -1625 7453 -1573
rect 7453 -1625 7478 -1573
rect 7509 -1625 7517 -1573
rect 7517 -1625 7565 -1573
rect 7596 -1625 7633 -1573
rect 7633 -1625 7645 -1573
rect 7645 -1625 7652 -1573
rect 7683 -1625 7697 -1573
rect 7697 -1625 7709 -1573
rect 7709 -1625 7739 -1573
rect 7770 -1625 7773 -1573
rect 7773 -1625 7825 -1573
rect 7825 -1625 7826 -1573
rect 5829 -1627 5885 -1625
rect 5921 -1627 5977 -1625
rect 6013 -1627 6069 -1625
rect 6105 -1627 6161 -1625
rect 6197 -1627 6253 -1625
rect 6289 -1627 6345 -1625
rect 6380 -1627 6436 -1625
rect 7247 -1627 7303 -1625
rect 7335 -1627 7391 -1625
rect 7422 -1627 7478 -1625
rect 7509 -1627 7565 -1625
rect 7596 -1627 7652 -1625
rect 7683 -1627 7739 -1625
rect 7770 -1627 7826 -1625
rect 6679 -1729 6735 -1727
rect 6766 -1729 6822 -1727
rect 6853 -1729 6909 -1727
rect 6679 -1781 6685 -1729
rect 6685 -1781 6735 -1729
rect 6766 -1781 6801 -1729
rect 6801 -1781 6813 -1729
rect 6813 -1781 6822 -1729
rect 6853 -1781 6865 -1729
rect 6865 -1781 6877 -1729
rect 6877 -1781 6909 -1729
rect 6679 -1783 6735 -1781
rect 6766 -1783 6822 -1781
rect 6853 -1783 6909 -1781
rect 5829 -1885 5885 -1883
rect 5921 -1885 5977 -1883
rect 6013 -1885 6069 -1883
rect 6105 -1885 6161 -1883
rect 6197 -1885 6253 -1883
rect 6289 -1885 6345 -1883
rect 6380 -1885 6436 -1883
rect 7247 -1885 7303 -1883
rect 7335 -1885 7391 -1883
rect 7422 -1885 7478 -1883
rect 7509 -1885 7565 -1883
rect 7596 -1885 7652 -1883
rect 7683 -1885 7739 -1883
rect 7770 -1885 7826 -1883
rect 5829 -1937 5846 -1885
rect 5846 -1937 5885 -1885
rect 5921 -1937 5963 -1885
rect 5963 -1937 5976 -1885
rect 5976 -1937 5977 -1885
rect 6013 -1937 6028 -1885
rect 6028 -1937 6041 -1885
rect 6041 -1937 6069 -1885
rect 6105 -1937 6106 -1885
rect 6106 -1937 6158 -1885
rect 6158 -1937 6161 -1885
rect 6197 -1937 6223 -1885
rect 6223 -1937 6236 -1885
rect 6236 -1937 6253 -1885
rect 6289 -1937 6301 -1885
rect 6301 -1937 6345 -1885
rect 6380 -1937 6417 -1885
rect 6417 -1937 6429 -1885
rect 6429 -1937 6436 -1885
rect 7247 -1937 7249 -1885
rect 7249 -1937 7261 -1885
rect 7261 -1937 7303 -1885
rect 7335 -1937 7377 -1885
rect 7377 -1937 7389 -1885
rect 7389 -1937 7391 -1885
rect 7422 -1937 7441 -1885
rect 7441 -1937 7453 -1885
rect 7453 -1937 7478 -1885
rect 7509 -1937 7517 -1885
rect 7517 -1937 7565 -1885
rect 7596 -1937 7633 -1885
rect 7633 -1937 7645 -1885
rect 7645 -1937 7652 -1885
rect 7683 -1937 7697 -1885
rect 7697 -1937 7709 -1885
rect 7709 -1937 7739 -1885
rect 7770 -1937 7773 -1885
rect 7773 -1937 7825 -1885
rect 7825 -1937 7826 -1885
rect 5829 -1939 5885 -1937
rect 5921 -1939 5977 -1937
rect 6013 -1939 6069 -1937
rect 6105 -1939 6161 -1937
rect 6197 -1939 6253 -1937
rect 6289 -1939 6345 -1937
rect 6380 -1939 6436 -1937
rect 7247 -1939 7303 -1937
rect 7335 -1939 7391 -1937
rect 7422 -1939 7478 -1937
rect 7509 -1939 7565 -1937
rect 7596 -1939 7652 -1937
rect 7683 -1939 7739 -1937
rect 7770 -1939 7826 -1937
rect 6535 -2742 6591 -2686
rect 6535 -2822 6591 -2766
<< metal3 >>
rect 6274 1452 6792 1562
tri 6792 1452 6902 1562 sw
rect 6274 1447 6902 1452
rect 6274 1427 6679 1447
tri 6587 1391 6623 1427 ne
rect 6623 1391 6679 1427
rect 6735 1391 6759 1447
rect 6815 1391 6839 1447
rect 6895 1440 6902 1447
tri 6902 1440 6914 1452 sw
rect 6895 1391 6914 1440
tri 6623 1365 6649 1391 ne
rect 6649 1365 6914 1391
tri 6649 1340 6674 1365 ne
rect 5814 1269 6445 1338
rect 5814 1213 5823 1269
rect 5879 1213 5904 1269
rect 5960 1213 5984 1269
rect 6040 1213 6064 1269
rect 6120 1213 6144 1269
rect 6200 1213 6224 1269
rect 6280 1213 6304 1269
rect 6360 1213 6384 1269
rect 6440 1213 6445 1269
rect 5814 957 6445 1213
rect 5814 901 5823 957
rect 5879 901 5904 957
rect 5960 901 5984 957
rect 6040 901 6064 957
rect 6120 901 6144 957
rect 6200 901 6224 957
rect 6280 901 6304 957
rect 6360 901 6384 957
rect 6440 901 6445 957
rect 5814 645 6445 901
rect 5814 589 5823 645
rect 5879 589 5904 645
rect 5960 589 5984 645
rect 6040 589 6064 645
rect 6120 589 6144 645
rect 6200 589 6224 645
rect 6280 589 6304 645
rect 6360 589 6384 645
rect 6440 589 6445 645
rect 6674 1309 6679 1365
rect 6735 1309 6759 1365
rect 6815 1309 6839 1365
rect 6895 1309 6914 1365
rect 6674 1113 6914 1309
rect 6674 1057 6683 1113
rect 6739 1057 6766 1113
rect 6822 1057 6849 1113
rect 6905 1057 6914 1113
rect 6674 801 6914 1057
rect 6674 745 6683 801
rect 6739 745 6766 801
rect 6822 745 6849 801
rect 6905 745 6914 801
rect 5814 -1259 6445 589
rect 5814 -1315 5829 -1259
rect 5885 -1315 5921 -1259
rect 5977 -1315 6013 -1259
rect 6069 -1315 6105 -1259
rect 6161 -1315 6197 -1259
rect 6253 -1315 6289 -1259
rect 6345 -1315 6380 -1259
rect 6436 -1315 6445 -1259
rect 5814 -1571 6445 -1315
rect 5814 -1627 5829 -1571
rect 5885 -1627 5921 -1571
rect 5977 -1627 6013 -1571
rect 6069 -1627 6105 -1571
rect 6161 -1627 6197 -1571
rect 6253 -1627 6289 -1571
rect 6345 -1627 6380 -1571
rect 6436 -1627 6445 -1571
rect 5814 -1883 6445 -1627
rect 5814 -1939 5829 -1883
rect 5885 -1939 5921 -1883
rect 5977 -1939 6013 -1883
rect 6069 -1939 6105 -1883
rect 6161 -1939 6197 -1883
rect 6253 -1939 6289 -1883
rect 6345 -1939 6380 -1883
rect 6436 -1939 6445 -1883
rect 5814 -1944 6445 -1939
rect 6530 634 6596 639
rect 6530 578 6535 634
rect 6591 578 6596 634
rect 6530 554 6596 578
rect 6530 498 6535 554
rect 6591 498 6596 554
rect 6530 -2686 6596 498
rect 6674 470 6914 745
rect 6674 414 6687 470
rect 6743 414 6767 470
rect 6823 414 6847 470
rect 6903 414 6914 470
rect 6674 388 6914 414
rect 6674 332 6687 388
rect 6743 332 6767 388
rect 6823 332 6847 388
rect 6903 332 6914 388
rect 6674 -1415 6914 332
rect 6674 -1471 6679 -1415
rect 6735 -1471 6766 -1415
rect 6822 -1471 6853 -1415
rect 6909 -1471 6914 -1415
rect 6674 -1727 6914 -1471
rect 6674 -1783 6679 -1727
rect 6735 -1783 6766 -1727
rect 6822 -1783 6853 -1727
rect 6909 -1783 6914 -1727
rect 6674 -1788 6914 -1783
rect 7242 1269 8048 1342
rect 7242 1213 7427 1269
rect 7483 1213 7507 1269
rect 7563 1213 7587 1269
rect 7643 1213 7667 1269
rect 7723 1213 7747 1269
rect 7803 1213 7827 1269
rect 7883 1213 7907 1269
rect 7963 1213 7987 1269
rect 8043 1213 8048 1269
rect 7242 957 8048 1213
rect 7242 901 7427 957
rect 7483 901 7520 957
rect 7576 901 7612 957
rect 7668 901 7704 957
rect 7760 901 7796 957
rect 7852 901 7888 957
rect 7944 901 7980 957
rect 8036 901 8048 957
rect 7242 645 8048 901
rect 10452 1269 10781 1859
rect 10452 1213 10461 1269
rect 10517 1213 10546 1269
rect 10602 1213 10631 1269
rect 10687 1213 10716 1269
rect 10772 1213 10781 1269
rect 10452 957 10781 1213
rect 10452 901 10461 957
rect 10517 901 10546 957
rect 10602 901 10631 957
rect 10687 901 10716 957
rect 10772 901 10781 957
rect 10452 803 10781 901
rect 7242 589 7427 645
rect 7483 589 7507 645
rect 7563 589 7587 645
rect 7643 589 7667 645
rect 7723 589 7747 645
rect 7803 589 7827 645
rect 7883 589 7907 645
rect 7963 589 7987 645
rect 8043 589 8048 645
rect 7242 535 8048 589
rect 7242 438 7951 535
tri 7951 438 8048 535 nw
rect 10452 645 10781 736
rect 10452 589 10461 645
rect 10517 589 10546 645
rect 10602 589 10631 645
rect 10687 589 10716 645
rect 10772 589 10781 645
rect 10452 438 10781 589
rect 7242 -1259 7879 438
tri 7879 366 7951 438 nw
rect 7242 -1315 7247 -1259
rect 7303 -1315 7335 -1259
rect 7391 -1315 7422 -1259
rect 7478 -1315 7509 -1259
rect 7565 -1315 7596 -1259
rect 7652 -1315 7683 -1259
rect 7739 -1315 7770 -1259
rect 7826 -1315 7879 -1259
rect 7242 -1571 7879 -1315
rect 7242 -1627 7247 -1571
rect 7303 -1627 7335 -1571
rect 7391 -1627 7422 -1571
rect 7478 -1627 7509 -1571
rect 7565 -1627 7596 -1571
rect 7652 -1627 7683 -1571
rect 7739 -1627 7770 -1571
rect 7826 -1627 7879 -1571
rect 7242 -1883 7879 -1627
rect 7242 -1939 7247 -1883
rect 7303 -1939 7335 -1883
rect 7391 -1939 7422 -1883
rect 7478 -1939 7509 -1883
rect 7565 -1939 7596 -1883
rect 7652 -1939 7683 -1883
rect 7739 -1939 7770 -1883
rect 7826 -1939 7879 -1883
rect 7242 -1944 7879 -1939
rect 6530 -2742 6535 -2686
rect 6591 -2742 6596 -2686
rect 6530 -2766 6596 -2742
rect 6530 -2822 6535 -2766
rect 6591 -2822 6596 -2766
rect 6530 -2831 6596 -2822
use sky130_fd_pr__nfet_01v8__example_55959141808516  sky130_fd_pr__nfet_01v8__example_55959141808516_1
timestamp 1633016201
transform 0 1 558 -1 0 1187
box -28 0 284 471
use sky130_fd_pr__nfet_01v8__example_55959141808516  sky130_fd_pr__nfet_01v8__example_55959141808516_0
timestamp 1633016201
transform 0 1 558 -1 0 745
box -28 0 284 471
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_1
timestamp 1633016201
transform 0 -1 -104 1 0 612
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1633016201
transform 0 -1 -104 -1 0 694
box 0 0 882 404
use sky130_fd_pr__nfet_01v8__example_55959141808523  sky130_fd_pr__nfet_01v8__example_55959141808523_0
timestamp 1633016201
transform 0 -1 9412 -1 0 1213
box -28 0 752 981
use sky130_fd_pr__nfet_01v8__example_55959141808523  sky130_fd_pr__nfet_01v8__example_55959141808523_1
timestamp 1633016201
transform 0 -1 6499 1 0 489
box -28 0 752 981
use sky130_fd_pr__nfet_01v8__example_55959141808522  sky130_fd_pr__nfet_01v8__example_55959141808522_0
timestamp 1633016201
transform 0 -1 11518 1 0 801
box -28 0 440 981
use sky130_fd_pr__nfet_01v8__example_55959141808522  sky130_fd_pr__nfet_01v8__example_55959141808522_1
timestamp 1633016201
transform 0 1 2393 1 0 801
box -28 0 440 981
use sky130_fd_pr__nfet_01v8__example_55959141808519  sky130_fd_pr__nfet_01v8__example_55959141808519_0
timestamp 1633016201
transform 0 1 2393 1 0 489
box -28 0 284 981
use sky130_fd_pr__nfet_01v8__example_55959141808519  sky130_fd_pr__nfet_01v8__example_55959141808519_1
timestamp 1633016201
transform 0 -1 11518 1 0 489
box -28 0 284 981
use sky130_fd_pr__pfet_01v8__example_55959141808514  sky130_fd_pr__pfet_01v8__example_55959141808514_0
timestamp 1633016201
transform 0 -1 7816 1 0 -1883
box -28 0 596 981
<< labels >>
flabel metal3 s 6530 461 6596 513 3 FreeSans 520 0 0 0 NG_AG_VPMP
port 1 nsew
flabel metal3 s 5819 -611 6441 -234 3 FreeSans 520 0 0 0 AG_HV
port 2 nsew
flabel metal3 s 10455 1022 10772 1149 3 FreeSans 520 0 0 0 PAD_HV_N2
port 3 nsew
flabel metal3 s 10458 533 10775 681 3 FreeSans 520 0 0 0 PAD_HV_N3
port 4 nsew
flabel metal1 s -474 635 -185 762 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal2 s 3130 1095 3459 1225 3 FreeSans 520 0 0 0 PAD_HV_N0
port 6 nsew
flabel metal2 s 3131 633 3458 687 3 FreeSans 520 0 0 0 PAD_HV_N1
port 7 nsew
flabel metal2 s 467 550 519 586 3 FreeSans 520 0 0 0 NMID_VDDA
port 8 nsew
flabel metal2 s 2364 256 2472 288 3 FreeSans 520 0 0 0 NG_PAD_VPMP
port 9 nsew
flabel metal2 s 5724 -1404 5773 -1296 3 FreeSans 520 0 0 0 PG_AG_VDDA
port 10 nsew
flabel comment s 7150 628 7150 628 0 FreeSans 440 90 0 0 CONDIODE
flabel comment s 488 404 488 404 0 FreeSans 400 90 0 0 NMID_VDDA
flabel comment s 2150 628 2150 628 0 FreeSans 440 90 0 0 CONDIODE
flabel comment s 1602 223 1602 223 0 FreeSans 280 0 0 0 MID1
flabel comment s 1800 1075 1800 1075 0 FreeSans 280 0 0 0 MID
flabel comment s 292 628 292 628 0 FreeSans 440 90 0 0 CONDIODE
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48314532
string GDS_START 48027864
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016076
<< checkpaint >>
rect -1260 -1349 1554 1795
<< nwell >>
rect 0 0 294 472
<< pmos >>
rect 89 36 119 436
rect 175 36 205 436
<< pdiff >>
rect 36 397 89 436
rect 36 363 44 397
rect 78 363 89 397
rect 36 325 89 363
rect 36 291 44 325
rect 78 291 89 325
rect 36 253 89 291
rect 36 219 44 253
rect 78 219 89 253
rect 36 181 89 219
rect 36 147 44 181
rect 78 147 89 181
rect 36 109 89 147
rect 36 75 44 109
rect 78 75 89 109
rect 36 36 89 75
rect 119 397 175 436
rect 119 363 130 397
rect 164 363 175 397
rect 119 325 175 363
rect 119 291 130 325
rect 164 291 175 325
rect 119 253 175 291
rect 119 219 130 253
rect 164 219 175 253
rect 119 181 175 219
rect 119 147 130 181
rect 164 147 175 181
rect 119 109 175 147
rect 119 75 130 109
rect 164 75 175 109
rect 119 36 175 75
rect 205 397 258 436
rect 205 363 216 397
rect 250 363 258 397
rect 205 325 258 363
rect 205 291 216 325
rect 250 291 258 325
rect 205 253 258 291
rect 205 219 216 253
rect 250 219 258 253
rect 205 181 258 219
rect 205 147 216 181
rect 250 147 258 181
rect 205 109 258 147
rect 205 75 216 109
rect 250 75 258 109
rect 205 36 258 75
<< pdiffc >>
rect 44 363 78 397
rect 44 291 78 325
rect 44 219 78 253
rect 44 147 78 181
rect 44 75 78 109
rect 130 363 164 397
rect 130 291 164 325
rect 130 219 164 253
rect 130 147 164 181
rect 130 75 164 109
rect 216 363 250 397
rect 216 291 250 325
rect 216 219 250 253
rect 216 147 250 181
rect 216 75 250 109
<< poly >>
rect 80 519 214 535
rect 80 485 96 519
rect 130 485 164 519
rect 198 485 214 519
rect 80 467 214 485
rect 89 462 205 467
rect 89 436 119 462
rect 175 436 205 462
rect 89 10 119 36
rect 175 10 205 36
<< polycont >>
rect 96 485 130 519
rect 164 485 198 519
<< locali >>
rect 80 519 214 535
rect 80 485 94 519
rect 130 485 164 519
rect 200 485 214 519
rect 80 467 214 485
rect 44 397 78 421
rect 44 325 78 363
rect 44 253 78 291
rect 44 181 78 219
rect 44 109 78 147
rect 44 47 78 75
rect 130 397 164 421
rect 130 325 164 363
rect 130 253 164 291
rect 130 181 164 219
rect 130 109 164 147
rect 130 51 164 75
rect 216 397 250 421
rect 216 325 250 363
rect 216 253 250 291
rect 216 181 250 219
rect 216 109 250 147
rect 216 51 250 75
<< viali >>
rect 94 485 96 519
rect 96 485 128 519
rect 166 485 198 519
rect 198 485 200 519
rect 44 363 78 397
rect 44 291 78 325
rect 44 219 78 253
rect 44 147 78 181
rect 44 75 78 109
rect 130 363 164 397
rect 130 291 164 325
rect 130 219 164 253
rect 130 147 164 181
rect 130 75 164 109
rect 216 363 250 397
rect 216 291 250 325
rect 216 219 250 253
rect 216 147 250 181
rect 216 75 250 109
<< metal1 >>
rect 82 519 212 531
rect 82 485 94 519
rect 128 485 166 519
rect 200 485 212 519
rect 82 473 212 485
rect 38 397 84 421
rect 38 363 44 397
rect 78 363 84 397
rect 38 325 84 363
rect 38 291 44 325
rect 78 291 84 325
rect 38 253 84 291
rect 38 219 44 253
rect 78 219 84 253
rect 38 181 84 219
rect 38 147 44 181
rect 78 147 84 181
rect 38 109 84 147
rect 38 75 44 109
rect 78 75 84 109
rect 38 -29 84 75
rect 121 410 173 421
rect 121 346 173 358
rect 121 291 130 294
rect 164 291 173 294
rect 121 253 173 291
rect 121 219 130 253
rect 164 219 173 253
rect 121 181 173 219
rect 121 147 130 181
rect 164 147 173 181
rect 121 109 173 147
rect 121 75 130 109
rect 164 75 173 109
rect 121 51 173 75
rect 210 397 256 421
rect 210 363 216 397
rect 250 363 256 397
rect 210 325 256 363
rect 210 291 216 325
rect 250 291 256 325
rect 210 253 256 291
rect 210 219 216 253
rect 250 219 256 253
rect 210 181 256 219
rect 210 147 216 181
rect 250 147 256 181
rect 210 109 256 147
rect 210 75 216 109
rect 250 75 256 109
rect 210 -29 256 75
rect 38 -89 256 -29
<< via1 >>
rect 121 397 173 410
rect 121 363 130 397
rect 130 363 164 397
rect 164 363 173 397
rect 121 358 173 363
rect 121 325 173 346
rect 121 294 130 325
rect 130 294 164 325
rect 164 294 173 325
<< metal2 >>
rect 121 410 173 416
rect 121 346 173 358
rect 121 288 173 294
<< labels >>
flabel metal2 s 121 288 173 416 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 82 473 212 531 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 38 -89 256 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel nwell s 74 464 78 471 0 FreeSans 400 0 0 0 BULK
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9181656
string GDS_START 9176656
string path 5.825 10.525 5.825 -2.225 
<< end >>

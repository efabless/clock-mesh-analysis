magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -2133 -4026 16575 33110
<< locali >>
rect 410 16553 502 16599
rect 1019 15138 1058 15172
rect 1092 15138 1131 15172
rect 1165 15138 1204 15172
rect 1238 15138 1277 15172
rect 1311 15138 1350 15172
rect 1384 15138 1423 15172
rect 1457 15138 1496 15172
rect 1530 15138 1569 15172
rect 1603 15138 1642 15172
rect 1676 15138 1715 15172
rect 1749 15138 1788 15172
rect 1822 15138 1861 15172
rect 1895 15138 1934 15172
rect 1968 15138 2007 15172
rect 2041 15138 2080 15172
rect 2114 15138 2153 15172
rect 2187 15138 2226 15172
rect 2260 15138 2299 15172
rect 2333 15138 2372 15172
rect 2406 15138 2445 15172
rect 2479 15138 2518 15172
rect 2552 15138 2591 15172
rect 2625 15138 2664 15172
rect 2698 15138 2737 15172
rect 2771 15138 2810 15172
rect 2844 15138 2883 15172
rect 2917 15138 2956 15172
rect 2990 15138 3029 15172
rect 3063 15138 3102 15172
rect 3136 15138 3175 15172
rect 3209 15138 3248 15172
rect 3282 15138 3321 15172
rect 3355 15138 3394 15172
rect 3428 15138 3467 15172
rect 3501 15138 3540 15172
rect 3574 15138 3613 15172
rect 3647 15138 3686 15172
rect 3720 15138 3759 15172
rect 3793 15138 3832 15172
rect 3866 15138 3905 15172
rect 3939 15138 3978 15172
rect 4012 15138 4051 15172
rect 4085 15138 4124 15172
rect 4158 15138 4197 15172
rect 4231 15138 4270 15172
rect 4304 15138 4343 15172
rect 4377 15138 4416 15172
rect 4450 15138 4489 15172
rect 4523 15138 4562 15172
rect 4596 15138 4635 15172
rect 4669 15138 4708 15172
rect 4742 15138 4781 15172
rect 4815 15138 4853 15172
rect 4887 15138 4925 15172
rect 4959 15138 4997 15172
rect 5031 15138 5069 15172
rect 5103 15138 5141 15172
rect 5175 15138 5213 15172
rect 5247 15138 5285 15172
rect 5319 15138 5357 15172
rect 5391 15138 5429 15172
rect 5463 15138 5501 15172
rect 5535 15138 5573 15172
rect 5607 15138 5645 15172
rect 5679 15138 5717 15172
rect 5751 15138 5789 15172
rect 5823 15138 5861 15172
rect 5895 15138 5933 15172
rect 5967 15138 6005 15172
rect 6039 15138 6077 15172
rect 6111 15138 6149 15172
rect 6183 15138 6221 15172
rect 6255 15138 6293 15172
rect 6327 15138 6365 15172
rect 6399 15138 6437 15172
rect 6471 15138 6509 15172
rect 6543 15138 6581 15172
rect 6615 15138 6653 15172
rect 6687 15138 6725 15172
rect 6759 15138 6797 15172
rect 6831 15138 6869 15172
rect 6903 15138 6941 15172
rect 6975 15138 7013 15172
rect 7047 15138 7085 15172
rect 7119 15138 7157 15172
rect 7191 15138 7229 15172
rect 162 2283 208 2362
rect 162 2249 168 2283
rect 202 2249 208 2283
rect 162 2211 208 2249
rect 162 2177 168 2211
rect 202 2177 208 2211
rect 162 2139 208 2177
rect 162 2105 168 2139
rect 202 2105 208 2139
rect 162 2067 208 2105
rect 162 2033 168 2067
rect 202 2033 208 2067
rect 162 1995 208 2033
rect 162 1961 168 1995
rect 202 1961 208 1995
rect 162 1923 208 1961
rect 162 1889 168 1923
rect 202 1889 208 1923
rect 162 1851 208 1889
rect 162 1817 168 1851
rect 202 1817 208 1851
rect 162 1779 208 1817
rect 162 1745 168 1779
rect 202 1745 208 1779
rect 162 1707 208 1745
rect 162 1673 168 1707
rect 202 1673 208 1707
rect 162 1635 208 1673
rect 162 1601 168 1635
rect 202 1601 208 1635
rect 162 1563 208 1601
rect 162 1529 168 1563
rect 202 1529 208 1563
rect 162 1491 208 1529
rect 162 1457 168 1491
rect 202 1457 208 1491
rect 162 1419 208 1457
rect 162 1385 168 1419
rect 202 1385 208 1419
rect 162 1347 208 1385
rect 162 1313 168 1347
rect 202 1313 208 1347
rect 162 1275 208 1313
rect 162 1241 168 1275
rect 202 1241 208 1275
rect 162 1203 208 1241
rect 162 1169 168 1203
rect 202 1169 208 1203
rect 162 1131 208 1169
rect 162 1097 168 1131
rect 202 1097 208 1131
rect 162 1059 208 1097
rect 10701 1064 10807 1606
rect 10999 1064 11105 1606
rect 162 1025 168 1059
rect 202 1025 208 1059
rect 162 987 208 1025
rect 162 953 168 987
rect 202 953 208 987
rect 162 915 208 953
rect 162 881 168 915
rect 202 881 208 915
rect 162 843 208 881
rect 162 809 168 843
rect 202 809 208 843
rect 162 771 208 809
rect 162 737 168 771
rect 202 737 208 771
rect 162 699 208 737
rect 162 665 168 699
rect 202 665 208 699
rect 162 627 208 665
rect 162 593 168 627
rect 202 593 208 627
rect 162 555 208 593
rect 162 521 168 555
rect 202 521 208 555
rect 162 483 208 521
rect 162 449 168 483
rect 202 449 208 483
rect 162 411 208 449
rect 162 377 168 411
rect 202 377 208 411
rect 162 339 208 377
rect 162 305 168 339
rect 202 305 208 339
rect 162 267 208 305
rect 162 233 168 267
rect 202 233 208 267
rect 162 195 208 233
rect 162 161 168 195
rect 202 161 208 195
rect 162 123 208 161
rect 162 89 168 123
rect 202 89 208 123
rect 162 51 208 89
rect 162 17 168 51
rect 202 17 208 51
rect 162 -21 208 17
rect 162 -55 168 -21
rect 202 -55 208 -21
rect 162 -93 208 -55
rect 162 -127 168 -93
rect 202 -127 208 -93
rect 162 -165 208 -127
rect 162 -199 168 -165
rect 202 -199 208 -165
rect 162 -237 208 -199
rect 162 -271 168 -237
rect 202 -271 208 -237
rect 162 -309 208 -271
rect 162 -343 168 -309
rect 202 -343 208 -309
rect 162 -381 208 -343
rect 162 -415 168 -381
rect 202 -387 12291 -381
rect 202 -415 293 -387
rect 162 -421 293 -415
rect 327 -421 365 -387
rect 399 -421 437 -387
rect 471 -421 509 -387
rect 543 -421 581 -387
rect 615 -421 653 -387
rect 687 -421 725 -387
rect 759 -421 797 -387
rect 831 -421 869 -387
rect 903 -421 941 -387
rect 975 -421 1013 -387
rect 1047 -421 1085 -387
rect 1119 -421 1157 -387
rect 1191 -421 1229 -387
rect 1263 -421 1301 -387
rect 1335 -421 1373 -387
rect 1407 -421 1445 -387
rect 1479 -421 1517 -387
rect 1551 -421 1589 -387
rect 1623 -421 1661 -387
rect 1695 -421 1733 -387
rect 1767 -421 1805 -387
rect 1839 -421 1877 -387
rect 1911 -421 1949 -387
rect 1983 -421 2021 -387
rect 2055 -421 2093 -387
rect 2127 -421 2165 -387
rect 2199 -421 2237 -387
rect 2271 -421 2309 -387
rect 2343 -421 2381 -387
rect 2415 -421 2453 -387
rect 2487 -421 2525 -387
rect 2559 -421 2597 -387
rect 2631 -421 2669 -387
rect 2703 -421 2741 -387
rect 2775 -421 2813 -387
rect 2847 -421 2885 -387
rect 2919 -421 2957 -387
rect 2991 -421 3029 -387
rect 3063 -421 3101 -387
rect 3135 -421 3173 -387
rect 3207 -421 3245 -387
rect 3279 -421 3317 -387
rect 3351 -421 3389 -387
rect 3423 -421 3461 -387
rect 3495 -421 3533 -387
rect 3567 -421 3605 -387
rect 3639 -421 3677 -387
rect 3711 -421 3749 -387
rect 3783 -421 3821 -387
rect 3855 -421 3893 -387
rect 3927 -421 3965 -387
rect 3999 -421 4037 -387
rect 4071 -421 4109 -387
rect 4143 -421 4181 -387
rect 4215 -421 4253 -387
rect 4287 -421 4325 -387
rect 4359 -421 4397 -387
rect 4431 -421 4469 -387
rect 4503 -421 4541 -387
rect 4575 -421 4613 -387
rect 4647 -421 4685 -387
rect 4719 -421 4757 -387
rect 4791 -421 4829 -387
rect 4863 -421 4901 -387
rect 4935 -421 4973 -387
rect 5007 -421 5045 -387
rect 5079 -421 5117 -387
rect 5151 -421 5189 -387
rect 5223 -421 5261 -387
rect 5295 -421 5333 -387
rect 5367 -421 5405 -387
rect 5439 -421 5477 -387
rect 5511 -421 5549 -387
rect 5583 -421 5621 -387
rect 5655 -421 5693 -387
rect 5727 -421 5765 -387
rect 5799 -421 5837 -387
rect 5871 -421 5909 -387
rect 5943 -421 5981 -387
rect 6015 -421 6053 -387
rect 6087 -421 6125 -387
rect 6159 -421 6197 -387
rect 6231 -421 6269 -387
rect 6303 -421 6341 -387
rect 6375 -421 6413 -387
rect 6447 -421 6485 -387
rect 6519 -421 6557 -387
rect 6591 -421 6629 -387
rect 6663 -421 6701 -387
rect 6735 -421 6773 -387
rect 6807 -421 6845 -387
rect 6879 -421 6917 -387
rect 6951 -421 6989 -387
rect 7023 -421 7061 -387
rect 7095 -421 7133 -387
rect 7167 -421 7205 -387
rect 7239 -421 7277 -387
rect 7311 -421 7349 -387
rect 7383 -421 7421 -387
rect 7455 -421 7493 -387
rect 7527 -421 7565 -387
rect 7599 -421 7637 -387
rect 7671 -421 7709 -387
rect 7743 -421 7781 -387
rect 7815 -421 7853 -387
rect 7887 -421 7925 -387
rect 7959 -421 7997 -387
rect 8031 -421 8069 -387
rect 8103 -421 8141 -387
rect 8175 -421 8213 -387
rect 8247 -421 8285 -387
rect 8319 -421 8357 -387
rect 8391 -421 8429 -387
rect 8463 -421 8501 -387
rect 8535 -421 8573 -387
rect 8607 -421 8645 -387
rect 8679 -421 8717 -387
rect 8751 -421 8789 -387
rect 8823 -421 8861 -387
rect 8895 -421 8933 -387
rect 8967 -421 9005 -387
rect 9039 -421 9077 -387
rect 9111 -421 9149 -387
rect 9183 -421 9221 -387
rect 9255 -421 9293 -387
rect 9327 -421 9365 -387
rect 9399 -421 9437 -387
rect 9471 -421 9509 -387
rect 9543 -421 9581 -387
rect 9615 -421 9653 -387
rect 9687 -421 9725 -387
rect 9759 -421 9797 -387
rect 9831 -421 9869 -387
rect 9903 -421 9941 -387
rect 9975 -421 10013 -387
rect 10047 -421 10085 -387
rect 10119 -421 10157 -387
rect 10191 -421 10229 -387
rect 10263 -421 10301 -387
rect 10335 -421 10373 -387
rect 10407 -421 10445 -387
rect 10479 -421 10517 -387
rect 10551 -421 10589 -387
rect 10623 -421 10661 -387
rect 10695 -421 10733 -387
rect 10767 -421 10805 -387
rect 10839 -421 10877 -387
rect 10911 -421 10949 -387
rect 10983 -421 11021 -387
rect 11055 -421 11093 -387
rect 11127 -421 11165 -387
rect 11199 -421 11237 -387
rect 11271 -421 11309 -387
rect 11343 -421 11381 -387
rect 11415 -421 11453 -387
rect 11487 -421 11525 -387
rect 11559 -421 11597 -387
rect 11631 -421 11669 -387
rect 11703 -421 11741 -387
rect 11775 -421 11813 -387
rect 11847 -421 11885 -387
rect 11919 -421 11957 -387
rect 11991 -421 12029 -387
rect 12063 -421 12101 -387
rect 12135 -421 12173 -387
rect 12207 -421 12245 -387
rect 12279 -421 12291 -387
rect 162 -427 12293 -421
rect 7986 -433 12293 -427
<< viali >>
rect 985 15138 1019 15172
rect 1058 15138 1092 15172
rect 1131 15138 1165 15172
rect 1204 15138 1238 15172
rect 1277 15138 1311 15172
rect 1350 15138 1384 15172
rect 1423 15138 1457 15172
rect 1496 15138 1530 15172
rect 1569 15138 1603 15172
rect 1642 15138 1676 15172
rect 1715 15138 1749 15172
rect 1788 15138 1822 15172
rect 1861 15138 1895 15172
rect 1934 15138 1968 15172
rect 2007 15138 2041 15172
rect 2080 15138 2114 15172
rect 2153 15138 2187 15172
rect 2226 15138 2260 15172
rect 2299 15138 2333 15172
rect 2372 15138 2406 15172
rect 2445 15138 2479 15172
rect 2518 15138 2552 15172
rect 2591 15138 2625 15172
rect 2664 15138 2698 15172
rect 2737 15138 2771 15172
rect 2810 15138 2844 15172
rect 2883 15138 2917 15172
rect 2956 15138 2990 15172
rect 3029 15138 3063 15172
rect 3102 15138 3136 15172
rect 3175 15138 3209 15172
rect 3248 15138 3282 15172
rect 3321 15138 3355 15172
rect 3394 15138 3428 15172
rect 3467 15138 3501 15172
rect 3540 15138 3574 15172
rect 3613 15138 3647 15172
rect 3686 15138 3720 15172
rect 3759 15138 3793 15172
rect 3832 15138 3866 15172
rect 3905 15138 3939 15172
rect 3978 15138 4012 15172
rect 4051 15138 4085 15172
rect 4124 15138 4158 15172
rect 4197 15138 4231 15172
rect 4270 15138 4304 15172
rect 4343 15138 4377 15172
rect 4416 15138 4450 15172
rect 4489 15138 4523 15172
rect 4562 15138 4596 15172
rect 4635 15138 4669 15172
rect 4708 15138 4742 15172
rect 4781 15138 4815 15172
rect 4853 15138 4887 15172
rect 4925 15138 4959 15172
rect 4997 15138 5031 15172
rect 5069 15138 5103 15172
rect 5141 15138 5175 15172
rect 5213 15138 5247 15172
rect 5285 15138 5319 15172
rect 5357 15138 5391 15172
rect 5429 15138 5463 15172
rect 5501 15138 5535 15172
rect 5573 15138 5607 15172
rect 5645 15138 5679 15172
rect 5717 15138 5751 15172
rect 5789 15138 5823 15172
rect 5861 15138 5895 15172
rect 5933 15138 5967 15172
rect 6005 15138 6039 15172
rect 6077 15138 6111 15172
rect 6149 15138 6183 15172
rect 6221 15138 6255 15172
rect 6293 15138 6327 15172
rect 6365 15138 6399 15172
rect 6437 15138 6471 15172
rect 6509 15138 6543 15172
rect 6581 15138 6615 15172
rect 6653 15138 6687 15172
rect 6725 15138 6759 15172
rect 6797 15138 6831 15172
rect 6869 15138 6903 15172
rect 6941 15138 6975 15172
rect 7013 15138 7047 15172
rect 7085 15138 7119 15172
rect 7157 15138 7191 15172
rect 7229 15138 7263 15172
rect 168 2249 202 2283
rect 168 2177 202 2211
rect 168 2105 202 2139
rect 168 2033 202 2067
rect 168 1961 202 1995
rect 168 1889 202 1923
rect 168 1817 202 1851
rect 168 1745 202 1779
rect 168 1673 202 1707
rect 168 1601 202 1635
rect 168 1529 202 1563
rect 168 1457 202 1491
rect 168 1385 202 1419
rect 168 1313 202 1347
rect 168 1241 202 1275
rect 168 1169 202 1203
rect 168 1097 202 1131
rect 168 1025 202 1059
rect 168 953 202 987
rect 168 881 202 915
rect 168 809 202 843
rect 168 737 202 771
rect 168 665 202 699
rect 168 593 202 627
rect 168 521 202 555
rect 168 449 202 483
rect 168 377 202 411
rect 168 305 202 339
rect 168 233 202 267
rect 168 161 202 195
rect 168 89 202 123
rect 168 17 202 51
rect 168 -55 202 -21
rect 168 -127 202 -93
rect 168 -199 202 -165
rect 168 -271 202 -237
rect 168 -343 202 -309
rect 168 -415 202 -381
rect 293 -421 327 -387
rect 365 -421 399 -387
rect 437 -421 471 -387
rect 509 -421 543 -387
rect 581 -421 615 -387
rect 653 -421 687 -387
rect 725 -421 759 -387
rect 797 -421 831 -387
rect 869 -421 903 -387
rect 941 -421 975 -387
rect 1013 -421 1047 -387
rect 1085 -421 1119 -387
rect 1157 -421 1191 -387
rect 1229 -421 1263 -387
rect 1301 -421 1335 -387
rect 1373 -421 1407 -387
rect 1445 -421 1479 -387
rect 1517 -421 1551 -387
rect 1589 -421 1623 -387
rect 1661 -421 1695 -387
rect 1733 -421 1767 -387
rect 1805 -421 1839 -387
rect 1877 -421 1911 -387
rect 1949 -421 1983 -387
rect 2021 -421 2055 -387
rect 2093 -421 2127 -387
rect 2165 -421 2199 -387
rect 2237 -421 2271 -387
rect 2309 -421 2343 -387
rect 2381 -421 2415 -387
rect 2453 -421 2487 -387
rect 2525 -421 2559 -387
rect 2597 -421 2631 -387
rect 2669 -421 2703 -387
rect 2741 -421 2775 -387
rect 2813 -421 2847 -387
rect 2885 -421 2919 -387
rect 2957 -421 2991 -387
rect 3029 -421 3063 -387
rect 3101 -421 3135 -387
rect 3173 -421 3207 -387
rect 3245 -421 3279 -387
rect 3317 -421 3351 -387
rect 3389 -421 3423 -387
rect 3461 -421 3495 -387
rect 3533 -421 3567 -387
rect 3605 -421 3639 -387
rect 3677 -421 3711 -387
rect 3749 -421 3783 -387
rect 3821 -421 3855 -387
rect 3893 -421 3927 -387
rect 3965 -421 3999 -387
rect 4037 -421 4071 -387
rect 4109 -421 4143 -387
rect 4181 -421 4215 -387
rect 4253 -421 4287 -387
rect 4325 -421 4359 -387
rect 4397 -421 4431 -387
rect 4469 -421 4503 -387
rect 4541 -421 4575 -387
rect 4613 -421 4647 -387
rect 4685 -421 4719 -387
rect 4757 -421 4791 -387
rect 4829 -421 4863 -387
rect 4901 -421 4935 -387
rect 4973 -421 5007 -387
rect 5045 -421 5079 -387
rect 5117 -421 5151 -387
rect 5189 -421 5223 -387
rect 5261 -421 5295 -387
rect 5333 -421 5367 -387
rect 5405 -421 5439 -387
rect 5477 -421 5511 -387
rect 5549 -421 5583 -387
rect 5621 -421 5655 -387
rect 5693 -421 5727 -387
rect 5765 -421 5799 -387
rect 5837 -421 5871 -387
rect 5909 -421 5943 -387
rect 5981 -421 6015 -387
rect 6053 -421 6087 -387
rect 6125 -421 6159 -387
rect 6197 -421 6231 -387
rect 6269 -421 6303 -387
rect 6341 -421 6375 -387
rect 6413 -421 6447 -387
rect 6485 -421 6519 -387
rect 6557 -421 6591 -387
rect 6629 -421 6663 -387
rect 6701 -421 6735 -387
rect 6773 -421 6807 -387
rect 6845 -421 6879 -387
rect 6917 -421 6951 -387
rect 6989 -421 7023 -387
rect 7061 -421 7095 -387
rect 7133 -421 7167 -387
rect 7205 -421 7239 -387
rect 7277 -421 7311 -387
rect 7349 -421 7383 -387
rect 7421 -421 7455 -387
rect 7493 -421 7527 -387
rect 7565 -421 7599 -387
rect 7637 -421 7671 -387
rect 7709 -421 7743 -387
rect 7781 -421 7815 -387
rect 7853 -421 7887 -387
rect 7925 -421 7959 -387
rect 7997 -421 8031 -387
rect 8069 -421 8103 -387
rect 8141 -421 8175 -387
rect 8213 -421 8247 -387
rect 8285 -421 8319 -387
rect 8357 -421 8391 -387
rect 8429 -421 8463 -387
rect 8501 -421 8535 -387
rect 8573 -421 8607 -387
rect 8645 -421 8679 -387
rect 8717 -421 8751 -387
rect 8789 -421 8823 -387
rect 8861 -421 8895 -387
rect 8933 -421 8967 -387
rect 9005 -421 9039 -387
rect 9077 -421 9111 -387
rect 9149 -421 9183 -387
rect 9221 -421 9255 -387
rect 9293 -421 9327 -387
rect 9365 -421 9399 -387
rect 9437 -421 9471 -387
rect 9509 -421 9543 -387
rect 9581 -421 9615 -387
rect 9653 -421 9687 -387
rect 9725 -421 9759 -387
rect 9797 -421 9831 -387
rect 9869 -421 9903 -387
rect 9941 -421 9975 -387
rect 10013 -421 10047 -387
rect 10085 -421 10119 -387
rect 10157 -421 10191 -387
rect 10229 -421 10263 -387
rect 10301 -421 10335 -387
rect 10373 -421 10407 -387
rect 10445 -421 10479 -387
rect 10517 -421 10551 -387
rect 10589 -421 10623 -387
rect 10661 -421 10695 -387
rect 10733 -421 10767 -387
rect 10805 -421 10839 -387
rect 10877 -421 10911 -387
rect 10949 -421 10983 -387
rect 11021 -421 11055 -387
rect 11093 -421 11127 -387
rect 11165 -421 11199 -387
rect 11237 -421 11271 -387
rect 11309 -421 11343 -387
rect 11381 -421 11415 -387
rect 11453 -421 11487 -387
rect 11525 -421 11559 -387
rect 11597 -421 11631 -387
rect 11669 -421 11703 -387
rect 11741 -421 11775 -387
rect 11813 -421 11847 -387
rect 11885 -421 11919 -387
rect 11957 -421 11991 -387
rect 12029 -421 12063 -387
rect 12101 -421 12135 -387
rect 12173 -421 12207 -387
rect 12245 -421 12279 -387
<< metal1 >>
rect 2627 23516 2680 23562
rect 2747 23518 3011 23629
tri 3011 23518 3122 23629 sw
rect 2747 23514 5881 23518
rect 2747 23499 5681 23514
tri 2957 23388 3068 23499 ne
rect 3068 23462 5681 23499
rect 5733 23462 5746 23514
rect 5798 23462 5810 23514
rect 5862 23462 5881 23514
rect 3068 23440 5881 23462
rect 3068 23388 5681 23440
rect 5733 23388 5746 23440
rect 5798 23388 5810 23440
rect 5862 23388 5881 23440
rect 13410 23185 13465 23518
rect 551 16163 1720 16308
rect 11900 15967 11932 16025
tri 6705 15951 6710 15956 se
tri 6709 15904 6710 15905 ne
rect 6710 15904 6716 15956
rect 6768 15904 6780 15956
rect 6832 15904 6838 15956
rect 4219 15407 5388 15552
rect 14264 15319 14340 15371
tri 7129 15290 7158 15319 sw
rect 7129 15238 7158 15290
tri 7158 15238 7210 15290 sw
rect 7483 15238 7489 15290
rect 7541 15238 7555 15290
rect 7607 15287 7613 15290
tri 7613 15287 7616 15290 sw
tri 14397 15287 14400 15290 se
rect 7607 15238 14400 15287
tri 14400 15238 14401 15239 nw
rect 7129 15230 7210 15238
tri 7210 15230 7218 15238 sw
rect 973 15208 7218 15230
tri 832 15172 868 15208 ne
rect 868 15185 7218 15208
rect 868 15172 2309 15185
rect 2361 15172 2375 15185
tri 868 15138 902 15172 ne
rect 902 15138 985 15172
rect 1019 15138 1058 15172
rect 1092 15138 1131 15172
rect 1165 15138 1204 15172
rect 1238 15138 1277 15172
rect 1311 15138 1350 15172
rect 1384 15138 1423 15172
rect 1457 15138 1496 15172
rect 1530 15138 1569 15172
rect 1603 15138 1642 15172
rect 1676 15138 1715 15172
rect 1749 15138 1788 15172
rect 1822 15138 1861 15172
rect 1895 15138 1934 15172
rect 1968 15138 2007 15172
rect 2041 15138 2080 15172
rect 2114 15138 2153 15172
rect 2187 15138 2226 15172
rect 2260 15138 2299 15172
rect 2361 15138 2372 15172
tri 902 15067 973 15138 ne
rect 973 15133 2309 15138
rect 2361 15133 2375 15138
rect 2427 15133 2441 15185
rect 2493 15133 2506 15185
rect 2558 15133 2571 15185
rect 2623 15172 2636 15185
rect 2688 15172 2701 15185
rect 2753 15172 2766 15185
rect 2818 15172 2831 15185
rect 2883 15172 2896 15185
rect 2948 15178 7218 15185
tri 7218 15178 7270 15230 sw
rect 2948 15172 7275 15178
rect 2625 15138 2636 15172
rect 2698 15138 2701 15172
rect 2948 15138 2956 15172
rect 2990 15138 3029 15172
rect 3063 15138 3102 15172
rect 3136 15138 3175 15172
rect 3209 15138 3248 15172
rect 3282 15138 3321 15172
rect 3355 15138 3394 15172
rect 3428 15138 3467 15172
rect 3501 15138 3540 15172
rect 3574 15138 3613 15172
rect 3647 15138 3686 15172
rect 3720 15138 3759 15172
rect 3793 15138 3832 15172
rect 3866 15138 3905 15172
rect 3939 15138 3978 15172
rect 4012 15138 4051 15172
rect 4085 15138 4124 15172
rect 4158 15138 4197 15172
rect 4231 15138 4270 15172
rect 4304 15138 4343 15172
rect 4377 15138 4416 15172
rect 4450 15138 4489 15172
rect 4523 15138 4562 15172
rect 4596 15138 4635 15172
rect 4669 15138 4708 15172
rect 4742 15138 4781 15172
rect 4815 15138 4853 15172
rect 4887 15138 4925 15172
rect 4959 15138 4997 15172
rect 5031 15138 5069 15172
rect 5103 15138 5141 15172
rect 5175 15138 5213 15172
rect 5247 15138 5285 15172
rect 5319 15138 5357 15172
rect 5391 15138 5429 15172
rect 5463 15138 5501 15172
rect 5535 15138 5573 15172
rect 5607 15138 5645 15172
rect 5679 15138 5717 15172
rect 5751 15138 5789 15172
rect 5823 15138 5861 15172
rect 5895 15138 5933 15172
rect 5967 15138 6005 15172
rect 6039 15138 6077 15172
rect 6111 15138 6149 15172
rect 6183 15138 6221 15172
rect 6255 15138 6293 15172
rect 6327 15138 6365 15172
rect 6399 15138 6437 15172
rect 6471 15138 6509 15172
rect 6543 15138 6581 15172
rect 6615 15138 6653 15172
rect 6687 15138 6725 15172
rect 6759 15138 6797 15172
rect 6831 15138 6869 15172
rect 6903 15138 6941 15172
rect 6975 15138 7013 15172
rect 7047 15138 7085 15172
rect 7119 15138 7157 15172
rect 7191 15138 7229 15172
rect 7263 15138 7275 15172
rect 2623 15133 2636 15138
rect 2688 15133 2701 15138
rect 2753 15133 2766 15138
rect 2818 15133 2831 15138
rect 2883 15133 2896 15138
rect 2948 15133 7275 15138
rect 973 15132 7275 15133
tri 7275 15132 7316 15173 sw
rect 973 15055 7316 15132
tri 7316 15055 7393 15132 sw
tri 4747 14860 4921 15034 ne
rect 5007 14860 5071 14959
tri 5071 14860 5170 14959 nw
tri 5007 14796 5071 14860 nw
rect 56 13979 570 14325
tri 14553 6235 14560 6242 se
rect 14560 6235 14566 6242
tri 11948 6190 11993 6235 se
rect 11993 6195 14566 6235
rect 11993 6190 12006 6195
tri 12006 6190 12011 6195 nw
tri 14555 6190 14560 6195 ne
rect 14560 6190 14566 6195
rect 14618 6190 14630 6242
rect 14682 6190 14688 6242
rect 14722 6238 14774 6244
tri 11935 6177 11948 6190 se
rect 11948 6177 11993 6190
tri 11993 6177 12006 6190 nw
tri 14717 6177 14722 6182 se
rect 14722 6177 14774 6186
tri 11914 6156 11935 6177 se
rect 11935 6156 11972 6177
tri 11972 6156 11993 6177 nw
tri 14696 6156 14717 6177 se
rect 14717 6174 14774 6177
rect 14717 6156 14722 6174
tri 11901 6143 11914 6156 se
rect 11914 6143 11956 6156
rect 6258 6140 6310 6143
tri 6310 6140 6313 6143 sw
tri 11898 6140 11901 6143 se
rect 11901 6140 11956 6143
tri 11956 6140 11972 6156 nw
tri 12021 6140 12037 6156 se
rect 12037 6140 14722 6156
rect 6258 6137 11928 6140
rect 6310 6112 11928 6137
tri 11928 6112 11956 6140 nw
tri 11993 6112 12021 6140 se
rect 12021 6122 14722 6140
rect 12021 6116 14774 6122
rect 14802 6157 14854 6163
rect 12021 6112 12037 6116
rect 6310 6100 6636 6112
tri 6636 6100 6648 6112 nw
tri 11981 6100 11993 6112 se
rect 11993 6100 12037 6112
rect 6310 6098 6343 6100
tri 6343 6098 6345 6100 nw
tri 11979 6098 11981 6100 se
rect 11981 6098 12037 6100
tri 12037 6098 12055 6116 nw
tri 14797 6098 14802 6103 se
rect 14802 6098 14854 6105
rect 6310 6085 6329 6098
rect 6258 6084 6329 6085
tri 6329 6084 6343 6098 nw
tri 11965 6084 11979 6098 se
rect 11979 6084 12023 6098
tri 12023 6084 12037 6098 nw
tri 14783 6084 14797 6098 se
rect 14797 6093 14854 6098
rect 14797 6084 14802 6093
rect 5832 5732 5899 6080
rect 6258 6073 6310 6084
tri 6310 6065 6329 6084 nw
rect 7388 6032 7394 6084
rect 7446 6032 7458 6084
rect 7510 6075 12014 6084
tri 12014 6075 12023 6084 nw
tri 14774 6075 14783 6084 se
rect 14783 6075 14802 6084
rect 7510 6072 12011 6075
tri 12011 6072 12014 6075 nw
tri 12066 6072 12069 6075 se
rect 12069 6072 14802 6075
rect 7510 6044 11983 6072
tri 11983 6044 12011 6072 nw
tri 12038 6044 12066 6072 se
rect 12066 6044 14802 6072
rect 7510 6032 7516 6044
tri 7516 6032 7528 6044 nw
tri 12029 6035 12038 6044 se
rect 12038 6041 14802 6044
rect 12038 6035 14854 6041
rect 14882 6074 14934 6080
tri 12026 6032 12029 6035 se
rect 12029 6032 12069 6035
rect 6258 6015 6310 6021
tri 12011 6017 12026 6032 se
rect 12026 6017 12069 6032
tri 12069 6017 12087 6035 nw
tri 12010 6016 12011 6017 se
rect 12011 6016 12056 6017
rect 8166 5964 8172 6016
rect 8224 5964 8236 6016
rect 8288 6004 8294 6016
tri 8294 6004 8306 6016 sw
tri 11998 6004 12010 6016 se
rect 12010 6004 12056 6016
tri 12056 6004 12069 6017 nw
tri 14870 6004 14882 6016 se
rect 14882 6010 14934 6022
rect 8288 5988 12040 6004
tri 12040 5988 12056 6004 nw
tri 14854 5988 14870 6004 se
rect 14870 5988 14882 6004
rect 8288 5975 12027 5988
tri 12027 5975 12040 5988 nw
tri 12069 5975 12082 5988 se
rect 12082 5975 14882 5988
rect 8288 5964 12016 5975
tri 12016 5964 12027 5975 nw
tri 12058 5964 12069 5975 se
rect 12069 5964 14882 5975
tri 12030 5936 12058 5964 se
rect 12058 5958 14882 5964
rect 12058 5952 14934 5958
rect 14962 5994 15014 6000
rect 12058 5948 14912 5952
tri 14912 5948 14916 5952 nw
rect 12058 5936 12083 5948
rect 9186 5884 9192 5936
rect 9244 5884 9256 5936
rect 9308 5931 9314 5936
tri 9314 5931 9319 5936 sw
tri 12025 5931 12030 5936 se
rect 12030 5931 12083 5936
tri 12083 5931 12100 5948 nw
tri 14953 5931 14962 5940 se
rect 14962 5931 15014 5942
rect 9308 5914 12066 5931
tri 12066 5914 12083 5931 nw
tri 14936 5914 14953 5931 se
rect 14953 5930 15014 5931
rect 14953 5914 14962 5930
rect 9308 5912 12064 5914
tri 12064 5912 12066 5914 nw
tri 14934 5912 14936 5914 se
rect 14936 5912 14962 5914
rect 9308 5891 12043 5912
tri 12043 5891 12064 5912 nw
tri 12085 5891 12106 5912 se
rect 12106 5891 14962 5912
rect 9308 5884 9314 5891
tri 9314 5884 9321 5891 nw
tri 12078 5884 12085 5891 se
rect 12085 5884 14962 5891
tri 12057 5863 12078 5884 se
rect 12078 5878 14962 5884
rect 12078 5872 15014 5878
rect 15042 5908 15094 5914
rect 12078 5863 12115 5872
tri 12115 5863 12124 5872 nw
rect 9967 5811 9973 5863
rect 10025 5811 10037 5863
rect 10089 5823 12075 5863
tri 12075 5823 12115 5863 nw
tri 15018 5830 15042 5854 se
rect 15042 5844 15094 5856
rect 10089 5811 10095 5823
tri 10095 5811 10107 5823 nw
rect 12123 5778 12129 5830
rect 12181 5778 12193 5830
rect 12245 5778 12251 5830
rect 12304 5778 12310 5830
rect 12362 5778 12374 5830
rect 12426 5826 12432 5830
tri 12432 5826 12436 5830 sw
tri 15014 5826 15018 5830 se
rect 15018 5826 15042 5830
rect 12426 5792 15042 5826
rect 12426 5786 15094 5792
rect 12426 5778 12432 5786
tri 12432 5778 12440 5786 nw
rect 7961 5722 7967 5774
rect 8019 5722 8031 5774
rect 8083 5734 11940 5774
rect 8083 5722 8089 5734
tri 8089 5722 8101 5734 nw
tri 11922 5722 11934 5734 ne
rect 11934 5722 11940 5734
rect 11992 5722 12004 5774
rect 12056 5722 12062 5774
rect 14751 5639 14886 5756
rect 14721 5357 14764 5395
rect 277 5087 317 5289
rect 12999 5017 13039 5219
rect 13072 5034 13239 5190
rect 14371 4633 14423 4639
tri 7307 4569 7359 4621 se
rect 7359 4569 7641 4621
rect 7693 4569 7705 4621
rect 7757 4569 7763 4621
tri 7285 4547 7307 4569 se
rect 7307 4547 7359 4569
tri 7359 4547 7381 4569 nw
rect 14371 4563 14423 4581
rect 14934 4574 15008 4609
tri 7243 4505 7285 4547 se
rect 7285 4505 7317 4547
tri 7317 4505 7359 4547 nw
rect 14371 4505 14423 4511
tri 7211 4473 7243 4505 se
rect 7243 4473 7285 4505
tri 7285 4473 7317 4505 nw
tri 7144 4406 7211 4473 se
rect 7211 4406 7218 4473
tri 7218 4406 7285 4473 nw
rect 5816 4354 5822 4406
rect 5874 4354 5886 4406
rect 5938 4354 7166 4406
tri 7166 4354 7218 4406 nw
rect 422 4168 462 4298
rect 12433 4188 12600 4285
rect 12797 4169 12837 4298
tri 12947 4169 12999 4221 se
rect 12999 4169 13136 4221
tri 12946 4168 12947 4169 se
rect 12947 4168 13136 4169
tri 12918 4140 12946 4168 se
rect 12946 4140 13136 4168
rect 185 3938 225 4140
rect 4046 4139 4349 4140
rect 4046 4087 4052 4139
rect 4104 4087 4132 4139
rect 4184 4087 4212 4139
rect 4264 4087 4291 4139
rect 4343 4087 4349 4139
rect 4046 4065 4349 4087
rect 4046 4013 4052 4065
rect 4104 4013 4132 4065
rect 4184 4013 4212 4065
rect 4264 4013 4291 4065
rect 4343 4013 4349 4065
rect 4046 3991 4349 4013
rect 4046 3939 4052 3991
rect 4104 3939 4132 3991
rect 4184 3939 4212 3991
rect 4264 3939 4291 3991
rect 4343 3939 4349 3991
rect 4046 3938 4349 3939
rect 12882 4019 13136 4140
rect 13148 4040 13459 4215
rect 12882 3938 13131 4019
tri 13131 3938 13212 4019 nw
rect 10259 3856 10265 3908
rect 10317 3856 10329 3908
rect 10381 3856 11619 3908
rect 11671 3856 11683 3908
rect 11735 3856 11741 3908
rect 4046 3683 4052 3735
rect 4104 3683 4132 3735
rect 4184 3683 4212 3735
rect 4264 3683 4291 3735
rect 4343 3683 4349 3735
rect 4046 3663 4349 3683
rect 4046 3611 4052 3663
rect 4104 3611 4132 3663
rect 4184 3611 4212 3663
rect 4264 3611 4291 3663
rect 4343 3611 4349 3663
tri 12194 3578 12195 3579 ne
rect 12195 3578 12244 3579
rect 5768 3521 5774 3573
rect 5826 3521 5838 3573
rect 5890 3521 7356 3573
rect 7408 3521 7420 3573
rect 7472 3521 7478 3573
rect 7537 3526 7543 3578
rect 7595 3526 7607 3578
rect 7659 3526 11609 3578
rect 11661 3526 11673 3578
rect 11725 3526 11731 3578
tri 12195 3529 12244 3578 ne
rect 14737 3488 14904 3644
rect 367 3209 409 3411
rect 8924 3209 8966 3411
tri 9994 3403 9997 3406 se
tri 9994 3354 9997 3357 ne
rect 9997 3354 10003 3406
rect 10055 3354 10067 3406
rect 10119 3354 10125 3406
tri 10125 3403 10128 3406 sw
tri 10125 3354 10128 3357 nw
rect 12437 3035 12489 3041
tri 12375 2965 12437 3027 se
rect 12437 2971 12489 2983
rect 11228 2913 11260 2965
rect 11312 2913 11324 2965
rect 11376 2919 12437 2965
rect 11376 2913 12489 2919
tri 12892 2913 12922 2943 se
tri 12864 2885 12892 2913 se
rect 12892 2885 12922 2913
rect 848 2683 890 2885
rect 4046 2884 4349 2885
rect 4046 2832 4052 2884
rect 4104 2832 4132 2884
rect 4184 2832 4212 2884
rect 4264 2832 4291 2884
rect 4343 2832 4349 2884
rect 4046 2810 4349 2832
rect 4046 2758 4052 2810
rect 4104 2758 4132 2810
rect 4184 2758 4212 2810
rect 4264 2758 4291 2810
rect 4343 2758 4349 2810
rect 4046 2736 4349 2758
rect 4046 2684 4052 2736
rect 4104 2684 4132 2736
rect 4184 2684 4212 2736
rect 4264 2684 4291 2736
rect 4343 2684 4349 2736
rect 4046 2683 4349 2684
rect 12531 2683 12933 2885
rect 14641 2790 14917 2796
rect 14641 2738 14642 2790
rect 14694 2738 14716 2790
rect 14768 2738 14790 2790
rect 14842 2738 14864 2790
rect 14916 2738 14917 2790
rect 14641 2722 14917 2738
rect 14594 2715 14917 2722
tri 12466 2522 12627 2683 ne
rect 12627 2522 12646 2683
rect 2587 2470 2593 2522
rect 2645 2470 2657 2522
rect 2709 2470 2715 2522
tri 12627 2503 12646 2522 ne
rect 14594 2663 14642 2715
rect 14694 2663 14716 2715
rect 14768 2663 14790 2715
rect 14842 2663 14864 2715
rect 14916 2663 14917 2715
rect 14594 2640 14917 2663
rect 14594 2588 14642 2640
rect 14694 2588 14716 2640
rect 14768 2588 14790 2640
rect 14842 2588 14864 2640
rect 14916 2588 14917 2640
rect 14594 2564 14917 2588
rect 14594 2512 14642 2564
rect 14694 2512 14716 2564
rect 14768 2512 14790 2564
rect 14842 2512 14864 2564
rect 14916 2512 14917 2564
rect 14594 2490 14917 2512
rect 14641 2488 14917 2490
rect 14641 2436 14642 2488
rect 14694 2436 14716 2488
rect 14768 2436 14790 2488
rect 14842 2436 14864 2488
rect 14916 2436 14917 2488
rect 14641 2430 14917 2436
rect 162 2283 208 2362
rect 162 2249 168 2283
rect 202 2249 208 2283
rect 162 2211 208 2249
rect 162 2177 168 2211
rect 202 2177 208 2211
rect 162 2139 208 2177
rect 1150 2158 1192 2288
rect 12031 2158 12096 2288
tri 12787 2194 12794 2201 se
rect 12794 2194 13325 2201
tri 12753 2160 12787 2194 se
rect 12787 2161 13325 2194
rect 12787 2160 12811 2161
tri 12811 2160 12812 2161 nw
tri 13210 2160 13211 2161 ne
rect 13211 2160 13325 2161
tri 13325 2160 13359 2194 sw
tri 12751 2158 12753 2160 se
rect 12753 2158 12794 2160
tri 12736 2143 12751 2158 se
rect 12751 2143 12794 2158
tri 12794 2143 12811 2160 nw
tri 13211 2143 13228 2160 ne
rect 13228 2143 13246 2160
rect 162 2105 168 2139
rect 202 2105 208 2139
rect 162 2067 208 2105
tri 12678 2085 12736 2143 se
tri 12736 2085 12794 2143 nw
tri 13228 2125 13246 2143 ne
rect 162 2033 168 2067
rect 202 2033 208 2067
rect 162 1995 208 2033
tri 12620 2027 12678 2085 se
tri 12678 2027 12736 2085 nw
rect 162 1961 168 1995
rect 202 1961 208 1995
tri 12571 1978 12620 2027 se
rect 162 1923 208 1961
rect 162 1889 168 1923
rect 202 1889 208 1923
rect 162 1851 208 1889
rect 162 1817 168 1851
rect 202 1817 208 1851
rect 10814 1972 10866 1978
tri 12562 1969 12571 1978 se
rect 12571 1969 12620 1978
tri 12620 1969 12678 2027 nw
rect 10814 1908 10866 1920
tri 12504 1911 12562 1969 se
tri 12562 1911 12620 1969 nw
tri 12500 1907 12504 1911 se
rect 12504 1907 12546 1911
tri 10866 1862 10892 1888 sw
rect 10866 1856 10980 1862
rect 10814 1855 10980 1856
tri 10980 1855 10987 1862 sw
rect 11149 1855 11155 1907
rect 11207 1855 11219 1907
rect 11271 1895 11277 1907
tri 11277 1895 11289 1907 sw
tri 12488 1895 12500 1907 se
rect 12500 1895 12546 1907
tri 12546 1895 12562 1911 nw
rect 11271 1855 12506 1895
tri 12506 1855 12546 1895 nw
rect 10814 1850 10987 1855
tri 10987 1850 10992 1855 sw
rect 10814 1827 10992 1850
tri 10992 1827 11015 1850 sw
rect 10814 1826 11015 1827
tri 11015 1826 11016 1827 sw
tri 11461 1826 11462 1827 se
rect 11462 1826 12580 1827
tri 12580 1826 12581 1827 sw
rect 10814 1824 11016 1826
rect 162 1779 208 1817
tri 10964 1813 10975 1824 ne
rect 10975 1813 11016 1824
tri 11016 1813 11029 1826 sw
tri 11448 1813 11461 1826 se
rect 11461 1813 12534 1826
tri 10975 1808 10980 1813 ne
rect 10980 1808 12534 1813
rect 162 1745 168 1779
rect 202 1745 208 1779
tri 10980 1774 11014 1808 ne
rect 11014 1788 12534 1808
rect 11014 1774 11486 1788
tri 11486 1774 11500 1788 nw
tri 12520 1774 12534 1788 ne
tri 10914 1746 10920 1752 sw
rect 162 1707 208 1745
rect 162 1673 168 1707
rect 202 1673 208 1707
rect 162 1635 208 1673
rect 162 1601 168 1635
rect 202 1601 208 1635
rect 162 1563 208 1601
rect 162 1529 168 1563
rect 202 1529 208 1563
rect 855 1542 897 1672
rect 12155 1542 12197 1672
rect 14737 1648 14904 1804
rect 162 1491 208 1529
rect 162 1457 168 1491
rect 202 1457 208 1491
rect 162 1419 208 1457
rect 162 1385 168 1419
rect 202 1385 208 1419
rect 162 1347 208 1385
rect 162 1313 168 1347
rect 202 1313 208 1347
tri 11827 1334 11833 1340 se
rect 162 1275 208 1313
rect 11833 1288 11839 1340
rect 11891 1288 11903 1340
rect 11955 1288 11961 1340
rect 162 1241 168 1275
rect 202 1241 208 1275
rect 162 1203 208 1241
rect -666 1182 -532 1188
rect -614 1130 -584 1182
rect -666 1105 -532 1130
rect -614 1053 -584 1105
rect -666 1027 -532 1053
rect -614 975 -584 1027
rect -666 969 -532 975
rect 162 1169 168 1203
rect 202 1169 208 1203
rect 162 1131 208 1169
rect 162 1097 168 1131
rect 202 1097 208 1131
rect 162 1059 208 1097
rect 162 1025 168 1059
rect 202 1025 208 1059
rect 857 1058 899 1260
rect 12059 1058 12101 1260
rect 12572 1192 12674 1198
rect 12624 1140 12674 1192
rect 12572 1126 12674 1140
rect 12624 1074 12674 1126
rect 12572 1068 12674 1074
rect 162 987 208 1025
rect 162 953 168 987
rect 202 953 208 987
rect 162 915 208 953
rect 162 881 168 915
rect 202 881 208 915
rect 162 843 208 881
rect 162 809 168 843
rect 202 809 208 843
rect 11151 842 11157 894
rect 11209 842 11221 894
rect 11273 888 12624 894
rect 11273 842 12572 888
rect 162 771 208 809
tri 12538 808 12572 842 ne
rect 12572 824 12624 836
rect 162 737 168 771
rect 202 737 208 771
rect 12572 766 12624 772
rect 162 734 208 737
rect 162 699 227 734
rect 162 665 168 699
rect 202 665 227 699
rect 162 627 227 665
rect 162 593 168 627
rect 202 593 227 627
rect 162 555 227 593
rect 162 521 168 555
rect 202 532 227 555
rect 4046 733 4349 734
rect 4046 681 4052 733
rect 4104 681 4132 733
rect 4184 681 4212 733
rect 4264 681 4291 733
rect 4343 681 4349 733
rect 4046 659 4349 681
rect 4046 607 4052 659
rect 4104 607 4132 659
rect 4184 607 4212 659
rect 4264 607 4291 659
rect 4343 607 4349 659
rect 4046 585 4349 607
rect 4046 533 4052 585
rect 4104 533 4132 585
rect 4184 533 4212 585
rect 4264 533 4291 585
rect 4343 533 4349 585
rect 4046 532 4349 533
rect 12370 653 12575 734
tri 12575 653 12656 734 sw
rect 12370 569 12634 653
rect 14641 648 14917 654
rect 14641 604 14642 648
tri 12370 532 12407 569 ne
rect 12407 532 12634 569
rect 202 521 208 532
rect 162 483 208 521
rect 162 449 168 483
rect 202 449 208 483
rect 162 411 208 449
tri 12407 424 12515 532 ne
rect 12515 424 12634 532
rect 162 377 168 411
rect 202 377 208 411
tri 5999 404 6002 407 se
rect 6002 404 6075 407
rect 162 339 208 377
rect 162 305 168 339
rect 202 305 208 339
rect 162 267 208 305
rect 5570 398 5622 404
tri 5622 378 5648 404 sw
tri 5973 378 5999 404 se
rect 5999 378 6075 404
rect 5622 372 5648 378
tri 5648 372 5654 378 sw
tri 5967 372 5973 378 se
rect 5973 372 6075 378
rect 5622 348 5654 372
tri 5654 348 5678 372 sw
tri 5943 348 5967 372 se
rect 5967 355 6075 372
rect 6127 355 6139 407
rect 6191 355 6197 407
tri 7759 372 7765 378 ne
rect 7765 372 7771 424
rect 7823 372 7835 424
rect 7887 372 7893 424
tri 12515 383 12556 424 ne
rect 12556 383 12634 424
rect 14594 596 14642 604
rect 14694 596 14716 648
rect 14768 596 14790 648
rect 14842 596 14864 648
rect 14916 596 14917 648
rect 14594 577 14917 596
rect 14594 525 14642 577
rect 14694 525 14716 577
rect 14768 525 14790 577
rect 14842 525 14864 577
rect 14916 525 14917 577
rect 14594 506 14917 525
rect 14594 454 14642 506
rect 14694 454 14716 506
rect 14768 454 14790 506
rect 14842 454 14864 506
rect 14916 454 14917 506
rect 14594 434 14917 454
rect 14594 382 14642 434
rect 14694 382 14716 434
rect 14768 382 14790 434
rect 14842 382 14864 434
rect 14916 382 14917 434
rect 14594 372 14917 382
rect 14641 362 14917 372
rect 5967 348 6017 355
tri 6017 348 6024 355 nw
rect 5622 346 5678 348
rect 5570 334 5678 346
rect 5622 333 5678 334
tri 5678 333 5693 348 sw
tri 5928 333 5943 348 se
rect 5943 333 6002 348
tri 6002 333 6017 348 nw
rect 5622 320 5693 333
tri 5693 320 5706 333 sw
tri 5915 320 5928 333 se
rect 5928 320 5989 333
tri 5989 320 6002 333 nw
rect 5622 312 5981 320
tri 5981 312 5989 320 nw
rect 5622 282 5945 312
rect 5570 276 5945 282
tri 5945 276 5981 312 nw
rect 162 233 168 267
rect 202 233 208 267
rect 8045 260 8051 312
rect 8103 260 8117 312
rect 8169 260 8175 312
rect 9203 260 9209 312
rect 9261 260 9275 312
rect 9327 260 9333 312
tri 10177 296 10183 302 ne
rect 10183 296 10189 348
rect 10241 296 10253 348
rect 10305 296 10311 348
rect 14641 310 14642 362
rect 14694 310 14716 362
rect 14768 310 14790 362
rect 14842 310 14864 362
rect 14916 310 14917 362
rect 14641 304 14917 310
rect 162 195 208 233
rect 162 161 168 195
rect 202 161 208 195
rect 162 123 208 161
rect 162 89 168 123
rect 202 89 208 123
rect 162 51 208 89
rect 162 17 168 51
rect 202 20 208 51
rect 202 17 222 20
rect 162 -21 222 17
rect 162 -55 168 -21
rect 202 -55 222 -21
rect 162 -93 222 -55
rect 162 -127 168 -93
rect 202 -126 222 -93
rect 1462 -32 1468 20
rect 1520 -32 1543 20
rect 1595 -32 1618 20
rect 1670 -32 1693 20
rect 1745 -32 1768 20
rect 1820 -32 1842 20
rect 1894 -32 1900 20
rect 1462 -74 1900 -32
rect 1462 -126 1468 -74
rect 1520 -126 1543 -74
rect 1595 -126 1618 -74
rect 1670 -126 1693 -74
rect 1745 -126 1768 -74
rect 1820 -126 1842 -74
rect 1894 -126 1900 -74
rect 4046 -32 4052 20
rect 4104 -32 4132 20
rect 4184 -32 4212 20
rect 4264 -32 4291 20
rect 4343 -32 4349 20
rect 4046 -74 4349 -32
rect 4046 -126 4052 -74
rect 4104 -126 4132 -74
rect 4184 -126 4212 -74
rect 4264 -126 4291 -74
rect 4343 -126 4349 -74
rect 12536 -126 12573 20
rect 202 -127 208 -126
rect 162 -165 208 -127
rect 162 -199 168 -165
rect 202 -199 208 -165
rect 162 -237 208 -199
rect 162 -271 168 -237
rect 202 -271 208 -237
rect 162 -309 208 -271
rect 162 -343 168 -309
rect 202 -343 208 -309
rect 162 -381 208 -343
tri 1651 -381 1654 -378 se
rect 1654 -381 1660 -378
rect 162 -415 168 -381
rect 202 -387 1660 -381
rect 1712 -387 1751 -378
rect 1803 -387 1842 -378
rect 1894 -381 1900 -378
tri 1900 -381 1903 -378 sw
tri 4043 -381 4046 -378 se
rect 4046 -381 4052 -378
rect 1894 -387 4052 -381
rect 4104 -387 4132 -378
rect 4184 -387 4212 -378
rect 4264 -387 4291 -378
rect 4343 -381 4349 -378
tri 4349 -381 4352 -378 sw
rect 4343 -387 12291 -381
rect 202 -415 293 -387
rect 162 -421 293 -415
rect 327 -421 365 -387
rect 399 -421 437 -387
rect 471 -421 509 -387
rect 543 -421 581 -387
rect 615 -421 653 -387
rect 687 -421 725 -387
rect 759 -421 797 -387
rect 831 -421 869 -387
rect 903 -421 941 -387
rect 975 -421 1013 -387
rect 1047 -421 1085 -387
rect 1119 -421 1157 -387
rect 1191 -421 1229 -387
rect 1263 -421 1301 -387
rect 1335 -421 1373 -387
rect 1407 -421 1445 -387
rect 1479 -421 1517 -387
rect 1551 -421 1589 -387
rect 1623 -421 1660 -387
rect 1712 -421 1733 -387
rect 1803 -421 1805 -387
rect 1839 -421 1842 -387
rect 1911 -421 1949 -387
rect 1983 -421 2021 -387
rect 2055 -421 2093 -387
rect 2127 -421 2165 -387
rect 2199 -421 2237 -387
rect 2271 -421 2309 -387
rect 2343 -421 2381 -387
rect 2415 -421 2453 -387
rect 2487 -421 2525 -387
rect 2559 -421 2597 -387
rect 2631 -421 2669 -387
rect 2703 -421 2741 -387
rect 2775 -421 2813 -387
rect 2847 -421 2885 -387
rect 2919 -421 2957 -387
rect 2991 -421 3029 -387
rect 3063 -421 3101 -387
rect 3135 -421 3173 -387
rect 3207 -421 3245 -387
rect 3279 -421 3317 -387
rect 3351 -421 3389 -387
rect 3423 -421 3461 -387
rect 3495 -421 3533 -387
rect 3567 -421 3605 -387
rect 3639 -421 3677 -387
rect 3711 -421 3749 -387
rect 3783 -421 3821 -387
rect 3855 -421 3893 -387
rect 3927 -421 3965 -387
rect 3999 -421 4037 -387
rect 4104 -421 4109 -387
rect 4287 -421 4291 -387
rect 4359 -421 4397 -387
rect 4431 -421 4469 -387
rect 4503 -421 4541 -387
rect 4575 -421 4613 -387
rect 4647 -421 4685 -387
rect 4719 -421 4757 -387
rect 4791 -421 4829 -387
rect 4863 -421 4901 -387
rect 4935 -421 4973 -387
rect 5007 -421 5045 -387
rect 5079 -421 5117 -387
rect 5151 -421 5189 -387
rect 5223 -421 5261 -387
rect 5295 -421 5333 -387
rect 5367 -421 5405 -387
rect 5439 -421 5477 -387
rect 5511 -421 5549 -387
rect 5583 -421 5621 -387
rect 5655 -421 5693 -387
rect 5727 -421 5765 -387
rect 5799 -421 5837 -387
rect 5871 -421 5909 -387
rect 5943 -421 5981 -387
rect 6015 -421 6053 -387
rect 6087 -421 6125 -387
rect 6159 -421 6197 -387
rect 6231 -421 6269 -387
rect 6303 -421 6341 -387
rect 6375 -421 6413 -387
rect 6447 -421 6485 -387
rect 6519 -421 6557 -387
rect 6591 -421 6629 -387
rect 6663 -421 6701 -387
rect 6735 -421 6773 -387
rect 6807 -421 6845 -387
rect 6879 -421 6917 -387
rect 6951 -421 6989 -387
rect 7023 -421 7061 -387
rect 7095 -421 7133 -387
rect 7167 -421 7205 -387
rect 7239 -421 7277 -387
rect 7311 -421 7349 -387
rect 7383 -421 7421 -387
rect 7455 -421 7493 -387
rect 7527 -421 7565 -387
rect 7599 -421 7637 -387
rect 7671 -421 7709 -387
rect 7743 -421 7781 -387
rect 7815 -421 7853 -387
rect 7887 -421 7925 -387
rect 7959 -421 7997 -387
rect 8031 -421 8069 -387
rect 8103 -421 8141 -387
rect 8175 -421 8213 -387
rect 8247 -421 8285 -387
rect 8319 -421 8357 -387
rect 8391 -421 8429 -387
rect 8463 -421 8501 -387
rect 8535 -421 8573 -387
rect 8607 -421 8645 -387
rect 8679 -421 8717 -387
rect 8751 -421 8789 -387
rect 8823 -421 8861 -387
rect 8895 -421 8933 -387
rect 8967 -421 9005 -387
rect 9039 -421 9077 -387
rect 9111 -421 9149 -387
rect 9183 -421 9221 -387
rect 9255 -421 9293 -387
rect 9327 -421 9365 -387
rect 9399 -421 9437 -387
rect 9471 -421 9509 -387
rect 9543 -421 9581 -387
rect 9615 -421 9653 -387
rect 9687 -421 9725 -387
rect 9759 -421 9797 -387
rect 9831 -421 9869 -387
rect 9903 -421 9941 -387
rect 9975 -421 10013 -387
rect 10047 -421 10085 -387
rect 10119 -421 10157 -387
rect 10191 -421 10229 -387
rect 10263 -421 10301 -387
rect 10335 -421 10373 -387
rect 10407 -421 10445 -387
rect 10479 -421 10517 -387
rect 10551 -421 10589 -387
rect 10623 -421 10661 -387
rect 10695 -421 10733 -387
rect 10767 -421 10805 -387
rect 10839 -421 10877 -387
rect 10911 -421 10949 -387
rect 10983 -421 11021 -387
rect 11055 -421 11093 -387
rect 11127 -421 11165 -387
rect 11199 -421 11237 -387
rect 11271 -421 11309 -387
rect 11343 -421 11381 -387
rect 11415 -421 11453 -387
rect 11487 -421 11525 -387
rect 11559 -421 11597 -387
rect 11631 -421 11669 -387
rect 11703 -421 11741 -387
rect 11775 -421 11813 -387
rect 11847 -421 11885 -387
rect 11919 -421 11957 -387
rect 11991 -421 12029 -387
rect 12063 -421 12101 -387
rect 12135 -421 12173 -387
rect 12207 -421 12245 -387
rect 12279 -421 12291 -387
rect 162 -427 1660 -421
tri 1651 -430 1654 -427 ne
rect 1654 -430 1660 -427
rect 1712 -430 1751 -421
rect 1803 -430 1842 -421
rect 1894 -427 4052 -421
rect 1894 -430 1900 -427
tri 1900 -430 1903 -427 nw
tri 4043 -430 4046 -427 ne
rect 4046 -430 4052 -427
rect 4104 -430 4132 -421
rect 4184 -430 4212 -421
rect 4264 -430 4291 -421
rect 4343 -427 12291 -421
rect 4343 -430 4349 -427
tri 4349 -430 4352 -427 nw
rect 10438 -515 10444 -463
rect 10496 -515 10508 -463
rect 10560 -515 12331 -463
rect 12383 -515 12395 -463
rect 12447 -515 12453 -463
rect 14737 -509 14904 -353
rect 10551 -595 10557 -543
rect 10609 -595 10621 -543
rect 10673 -595 12331 -543
rect 12383 -595 12395 -543
rect 12447 -595 12453 -543
rect 2853 -2686 2859 -2634
rect 2911 -2686 2923 -2634
rect 2975 -2686 2981 -2634
rect 11464 -2766 11470 -2714
rect 11522 -2766 11534 -2714
rect 11586 -2766 11592 -2714
<< via1 >>
rect 5681 23462 5733 23514
rect 5746 23462 5798 23514
rect 5810 23462 5862 23514
rect 5681 23388 5733 23440
rect 5746 23388 5798 23440
rect 5810 23388 5862 23440
rect 6716 15904 6768 15956
rect 6780 15904 6832 15956
rect 7489 15238 7541 15290
rect 7555 15238 7607 15290
rect 2309 15172 2361 15185
rect 2375 15172 2427 15185
rect 2309 15138 2333 15172
rect 2333 15138 2361 15172
rect 2375 15138 2406 15172
rect 2406 15138 2427 15172
rect 2309 15133 2361 15138
rect 2375 15133 2427 15138
rect 2441 15172 2493 15185
rect 2441 15138 2445 15172
rect 2445 15138 2479 15172
rect 2479 15138 2493 15172
rect 2441 15133 2493 15138
rect 2506 15172 2558 15185
rect 2506 15138 2518 15172
rect 2518 15138 2552 15172
rect 2552 15138 2558 15172
rect 2506 15133 2558 15138
rect 2571 15172 2623 15185
rect 2636 15172 2688 15185
rect 2701 15172 2753 15185
rect 2766 15172 2818 15185
rect 2831 15172 2883 15185
rect 2896 15172 2948 15185
rect 2571 15138 2591 15172
rect 2591 15138 2623 15172
rect 2636 15138 2664 15172
rect 2664 15138 2688 15172
rect 2701 15138 2737 15172
rect 2737 15138 2753 15172
rect 2766 15138 2771 15172
rect 2771 15138 2810 15172
rect 2810 15138 2818 15172
rect 2831 15138 2844 15172
rect 2844 15138 2883 15172
rect 2896 15138 2917 15172
rect 2917 15138 2948 15172
rect 2571 15133 2623 15138
rect 2636 15133 2688 15138
rect 2701 15133 2753 15138
rect 2766 15133 2818 15138
rect 2831 15133 2883 15138
rect 2896 15133 2948 15138
rect 14566 6190 14618 6242
rect 14630 6190 14682 6242
rect 14722 6186 14774 6238
rect 6258 6085 6310 6137
rect 14722 6122 14774 6174
rect 14802 6105 14854 6157
rect 6258 6021 6310 6073
rect 7394 6032 7446 6084
rect 7458 6032 7510 6084
rect 14802 6041 14854 6093
rect 14882 6022 14934 6074
rect 8172 5964 8224 6016
rect 8236 5964 8288 6016
rect 14882 5958 14934 6010
rect 9192 5884 9244 5936
rect 9256 5884 9308 5936
rect 14962 5942 15014 5994
rect 14962 5878 15014 5930
rect 9973 5811 10025 5863
rect 10037 5811 10089 5863
rect 15042 5856 15094 5908
rect 12129 5778 12181 5830
rect 12193 5778 12245 5830
rect 12310 5778 12362 5830
rect 12374 5778 12426 5830
rect 15042 5792 15094 5844
rect 7967 5722 8019 5774
rect 8031 5722 8083 5774
rect 11940 5722 11992 5774
rect 12004 5722 12056 5774
rect 7641 4569 7693 4621
rect 7705 4569 7757 4621
rect 14371 4581 14423 4633
rect 14371 4511 14423 4563
rect 5822 4354 5874 4406
rect 5886 4354 5938 4406
rect 4052 4087 4104 4139
rect 4132 4087 4184 4139
rect 4212 4087 4264 4139
rect 4291 4087 4343 4139
rect 4052 4013 4104 4065
rect 4132 4013 4184 4065
rect 4212 4013 4264 4065
rect 4291 4013 4343 4065
rect 4052 3939 4104 3991
rect 4132 3939 4184 3991
rect 4212 3939 4264 3991
rect 4291 3939 4343 3991
rect 10265 3856 10317 3908
rect 10329 3856 10381 3908
rect 11619 3856 11671 3908
rect 11683 3856 11735 3908
rect 4052 3683 4104 3735
rect 4132 3683 4184 3735
rect 4212 3683 4264 3735
rect 4291 3683 4343 3735
rect 4052 3611 4104 3663
rect 4132 3611 4184 3663
rect 4212 3611 4264 3663
rect 4291 3611 4343 3663
rect 5774 3521 5826 3573
rect 5838 3521 5890 3573
rect 7356 3521 7408 3573
rect 7420 3521 7472 3573
rect 7543 3526 7595 3578
rect 7607 3526 7659 3578
rect 11609 3526 11661 3578
rect 11673 3526 11725 3578
rect 10003 3354 10055 3406
rect 10067 3354 10119 3406
rect 12437 2983 12489 3035
rect 11260 2913 11312 2965
rect 11324 2913 11376 2965
rect 12437 2919 12489 2971
rect 4052 2832 4104 2884
rect 4132 2832 4184 2884
rect 4212 2832 4264 2884
rect 4291 2832 4343 2884
rect 4052 2758 4104 2810
rect 4132 2758 4184 2810
rect 4212 2758 4264 2810
rect 4291 2758 4343 2810
rect 4052 2684 4104 2736
rect 4132 2684 4184 2736
rect 4212 2684 4264 2736
rect 4291 2684 4343 2736
rect 14642 2738 14694 2790
rect 14716 2738 14768 2790
rect 14790 2738 14842 2790
rect 14864 2738 14916 2790
rect 2593 2470 2645 2522
rect 2657 2470 2709 2522
rect 14642 2663 14694 2715
rect 14716 2663 14768 2715
rect 14790 2663 14842 2715
rect 14864 2663 14916 2715
rect 14642 2588 14694 2640
rect 14716 2588 14768 2640
rect 14790 2588 14842 2640
rect 14864 2588 14916 2640
rect 14642 2512 14694 2564
rect 14716 2512 14768 2564
rect 14790 2512 14842 2564
rect 14864 2512 14916 2564
rect 14642 2436 14694 2488
rect 14716 2436 14768 2488
rect 14790 2436 14842 2488
rect 14864 2436 14916 2488
rect 10814 1920 10866 1972
rect 10814 1856 10866 1908
rect 11155 1855 11207 1907
rect 11219 1855 11271 1907
rect 11839 1288 11891 1340
rect 11903 1288 11955 1340
rect -666 1130 -614 1182
rect -584 1130 -532 1182
rect -666 1053 -614 1105
rect -584 1053 -532 1105
rect -666 975 -614 1027
rect -584 975 -532 1027
rect 12572 1140 12624 1192
rect 12572 1074 12624 1126
rect 11157 842 11209 894
rect 11221 842 11273 894
rect 12572 836 12624 888
rect 12572 772 12624 824
rect 4052 681 4104 733
rect 4132 681 4184 733
rect 4212 681 4264 733
rect 4291 681 4343 733
rect 4052 607 4104 659
rect 4132 607 4184 659
rect 4212 607 4264 659
rect 4291 607 4343 659
rect 4052 533 4104 585
rect 4132 533 4184 585
rect 4212 533 4264 585
rect 4291 533 4343 585
rect 5570 346 5622 398
rect 6075 355 6127 407
rect 6139 355 6191 407
rect 7771 372 7823 424
rect 7835 372 7887 424
rect 14642 596 14694 648
rect 14716 596 14768 648
rect 14790 596 14842 648
rect 14864 596 14916 648
rect 14642 525 14694 577
rect 14716 525 14768 577
rect 14790 525 14842 577
rect 14864 525 14916 577
rect 14642 454 14694 506
rect 14716 454 14768 506
rect 14790 454 14842 506
rect 14864 454 14916 506
rect 14642 382 14694 434
rect 14716 382 14768 434
rect 14790 382 14842 434
rect 14864 382 14916 434
rect 5570 282 5622 334
rect 8051 260 8103 312
rect 8117 260 8169 312
rect 9209 260 9261 312
rect 9275 260 9327 312
rect 10189 296 10241 348
rect 10253 296 10305 348
rect 14642 310 14694 362
rect 14716 310 14768 362
rect 14790 310 14842 362
rect 14864 310 14916 362
rect 1468 -32 1520 20
rect 1543 -32 1595 20
rect 1618 -32 1670 20
rect 1693 -32 1745 20
rect 1768 -32 1820 20
rect 1842 -32 1894 20
rect 1468 -126 1520 -74
rect 1543 -126 1595 -74
rect 1618 -126 1670 -74
rect 1693 -126 1745 -74
rect 1768 -126 1820 -74
rect 1842 -126 1894 -74
rect 4052 -32 4104 20
rect 4132 -32 4184 20
rect 4212 -32 4264 20
rect 4291 -32 4343 20
rect 4052 -126 4104 -74
rect 4132 -126 4184 -74
rect 4212 -126 4264 -74
rect 4291 -126 4343 -74
rect 1660 -387 1712 -378
rect 1751 -387 1803 -378
rect 1842 -387 1894 -378
rect 4052 -387 4104 -378
rect 4132 -387 4184 -378
rect 4212 -387 4264 -378
rect 4291 -387 4343 -378
rect 1660 -421 1661 -387
rect 1661 -421 1695 -387
rect 1695 -421 1712 -387
rect 1751 -421 1767 -387
rect 1767 -421 1803 -387
rect 1842 -421 1877 -387
rect 1877 -421 1894 -387
rect 4052 -421 4071 -387
rect 4071 -421 4104 -387
rect 4132 -421 4143 -387
rect 4143 -421 4181 -387
rect 4181 -421 4184 -387
rect 4212 -421 4215 -387
rect 4215 -421 4253 -387
rect 4253 -421 4264 -387
rect 4291 -421 4325 -387
rect 4325 -421 4343 -387
rect 1660 -430 1712 -421
rect 1751 -430 1803 -421
rect 1842 -430 1894 -421
rect 4052 -430 4104 -421
rect 4132 -430 4184 -421
rect 4212 -430 4264 -421
rect 4291 -430 4343 -421
rect 10444 -515 10496 -463
rect 10508 -515 10560 -463
rect 12331 -515 12383 -463
rect 12395 -515 12447 -463
rect 10557 -595 10609 -543
rect 10621 -595 10673 -543
rect 12331 -595 12383 -543
rect 12395 -595 12447 -543
rect 2859 -2686 2911 -2634
rect 2923 -2686 2975 -2634
rect 11470 -2766 11522 -2714
rect 11534 -2766 11586 -2714
<< metal2 >>
rect 3381 28647 3571 28656
rect 3437 28591 3515 28647
rect 3381 28565 3571 28591
rect 3437 28509 3515 28565
rect 3381 28483 3571 28509
rect 3437 28427 3515 28483
rect 3381 28401 3571 28427
rect 3437 28345 3515 28401
rect 3381 28319 3571 28345
rect 3437 28263 3515 28319
rect 3381 28237 3571 28263
rect 3437 28181 3515 28237
rect 3381 28155 3571 28181
rect 3437 28099 3515 28155
rect 3381 28073 3571 28099
rect 3437 28017 3515 28073
rect 3381 27991 3571 28017
rect 3437 27935 3515 27991
rect 3381 27909 3571 27935
rect 3437 27853 3515 27909
rect 3381 27827 3571 27853
rect 4626 27838 7525 28365
rect 3437 27771 3515 27827
rect 3381 27745 3571 27771
rect 3437 27689 3515 27745
rect 3381 27662 3571 27689
rect 3437 27606 3515 27662
rect 3381 27579 3571 27606
rect 3437 27523 3515 27579
rect 3381 27514 3571 27523
rect 11216 26085 12757 27178
rect 5668 23642 5868 23651
rect 5724 23586 5812 23642
rect 5668 23548 5868 23586
rect 5724 23514 5812 23548
rect 5668 23462 5681 23492
rect 5733 23462 5746 23514
rect 5798 23462 5810 23514
rect 5862 23462 5868 23492
rect 5668 23453 5868 23462
rect 5724 23440 5812 23453
rect 5668 23388 5681 23397
rect 5733 23388 5746 23440
rect 5798 23388 5810 23440
rect 5862 23388 5868 23397
rect 11216 19247 12757 20340
rect 13427 17780 14596 18850
rect 6710 15904 6716 15956
rect 6768 15904 6780 15956
rect 6832 15951 6838 15956
tri 6838 15951 6843 15956 sw
rect 6832 15905 7543 15951
rect 6832 15904 6838 15905
tri 6838 15904 6839 15905 nw
tri 7413 15904 7414 15905 ne
rect 7414 15904 7543 15905
tri 7543 15904 7590 15951 sw
tri 7414 15881 7437 15904 ne
rect 7437 15881 7590 15904
tri 7590 15881 7613 15904 sw
tri 7437 15835 7483 15881 ne
rect 7483 15290 7613 15881
rect 14635 15523 14768 15563
rect 14635 15511 14636 15523
tri 14636 15511 14648 15523 nw
tri 14702 15511 14714 15523 ne
rect 14714 15511 14768 15523
tri 14714 15497 14728 15511 ne
tri 14626 15401 14651 15426 ne
rect 7483 15238 7489 15290
rect 7541 15238 7555 15290
rect 7607 15238 7613 15290
tri 14459 15238 14460 15239 ne
rect 14460 15238 14528 15239
tri 14460 15220 14478 15238 ne
rect 14478 15220 14528 15238
tri 2027 15208 2039 15220 ne
rect 2039 15208 2963 15220
tri 14478 15208 14490 15220 ne
tri 2039 15185 2062 15208 ne
rect 2062 15185 2963 15208
tri 2062 15158 2089 15185 ne
rect 2089 15158 2309 15185
tri 2089 15133 2114 15158 ne
rect 2114 15133 2309 15158
rect 2361 15133 2375 15185
rect 2427 15133 2441 15185
rect 2493 15133 2506 15185
rect 2558 15133 2571 15185
rect 2623 15133 2636 15185
rect 2688 15133 2701 15185
rect 2753 15133 2766 15185
rect 2818 15133 2831 15185
rect 2883 15133 2896 15185
rect 2948 15133 2963 15185
tri 2114 15095 2152 15133 ne
rect 2152 15095 2963 15133
tri 14345 15095 14408 15158 ne
tri 2152 15046 2201 15095 ne
rect 2201 15046 2963 15095
tri 14387 6716 14408 6737 se
rect 14408 6719 14448 15158
rect 14408 6716 14445 6719
tri 14445 6716 14448 6719 nw
tri 14350 6679 14387 6716 se
rect 14387 6679 14408 6716
tri 14408 6679 14445 6716 nw
tri 14453 6679 14490 6716 se
rect 14490 6700 14528 15220
tri 14333 6662 14350 6679 se
rect 14350 6662 14391 6679
tri 14391 6662 14408 6679 nw
tri 14436 6662 14453 6679 se
rect 14453 6662 14490 6679
tri 14490 6662 14528 6700 nw
tri 14292 6621 14333 6662 se
rect 14333 6634 14363 6662
tri 14363 6634 14391 6662 nw
tri 14408 6634 14436 6662 se
rect 14333 6621 14350 6634
tri 14350 6621 14363 6634 nw
tri 14395 6621 14408 6634 se
rect 14408 6621 14436 6634
tri 14279 6608 14292 6621 se
rect 14292 6608 14337 6621
tri 14337 6608 14350 6621 nw
tri 14382 6608 14395 6621 se
rect 14395 6608 14436 6621
tri 14436 6608 14490 6662 nw
tri 14272 6601 14279 6608 se
rect 14279 6601 14330 6608
tri 14330 6601 14337 6608 nw
tri 14375 6601 14382 6608 se
rect 14382 6601 14408 6608
rect 3251 6108 3297 6154
rect 3724 6115 3776 6154
rect 6258 6137 6310 6143
rect 6258 6073 6310 6085
tri 14263 6084 14272 6093 se
rect 14272 6084 14312 6601
tri 14312 6583 14330 6601 nw
tri 14357 6583 14375 6601 se
rect 14375 6583 14408 6601
tri 4935 4358 4958 4381 ne
rect 4958 4358 5043 4381
tri 5043 4358 5066 4381 nw
rect 4958 4354 5039 4358
tri 5039 4354 5043 4358 nw
rect 5816 4354 5822 4406
rect 5874 4354 5886 4406
rect 5938 4354 5944 4406
rect 4046 4139 4349 4140
rect 4046 4087 4052 4139
rect 4104 4087 4132 4139
rect 4184 4087 4212 4139
rect 4264 4087 4291 4139
rect 4343 4087 4349 4139
rect 4046 4065 4349 4087
rect 4046 4013 4052 4065
rect 4104 4013 4132 4065
rect 4184 4013 4212 4065
rect 4264 4013 4291 4065
rect 4343 4013 4349 4065
rect 4046 3991 4349 4013
rect 4046 3939 4052 3991
rect 4104 3939 4132 3991
rect 4184 3939 4212 3991
rect 4264 3939 4291 3991
rect 4343 3939 4349 3991
rect 4046 3735 4349 3939
rect 4046 3683 4052 3735
rect 4104 3683 4132 3735
rect 4184 3683 4212 3735
rect 4264 3683 4291 3735
rect 4343 3683 4349 3735
rect 4046 3663 4349 3683
rect 4046 3611 4052 3663
rect 4104 3611 4132 3663
rect 4184 3611 4212 3663
rect 4264 3611 4291 3663
rect 4343 3611 4349 3663
rect 4046 2884 4349 3611
rect 4046 2832 4052 2884
rect 4104 2832 4132 2884
rect 4184 2832 4212 2884
rect 4264 2832 4291 2884
rect 4343 2832 4349 2884
rect 4046 2810 4349 2832
rect 4046 2758 4052 2810
rect 4104 2758 4132 2810
rect 4184 2758 4212 2810
rect 4264 2758 4291 2810
rect 4343 2758 4349 2810
rect 4046 2736 4349 2758
rect 4046 2684 4052 2736
rect 4104 2684 4132 2736
rect 4184 2684 4212 2736
rect 4264 2684 4291 2736
rect 4343 2684 4349 2736
rect 2587 2470 2593 2522
rect 2645 2470 2657 2522
rect 2709 2470 2715 2522
rect 2587 2436 2653 2470
tri 2653 2436 2687 2470 nw
rect -666 1182 -532 1188
rect -614 1130 -584 1182
rect -666 1105 -532 1130
rect -614 1053 -584 1105
rect -666 1027 -532 1053
rect -614 975 -584 1027
rect -666 539 -532 975
tri 1428 20 1518 110 sw
rect 1428 -32 1468 20
rect 1520 -32 1543 20
rect 1595 -32 1618 20
rect 1670 -32 1693 20
rect 1745 -32 1768 20
rect 1820 -32 1842 20
rect 1894 -32 1900 20
rect 1428 -74 1900 -32
rect 1428 -126 1468 -74
rect 1520 -126 1543 -74
rect 1595 -126 1618 -74
rect 1670 -126 1693 -74
rect 1745 -126 1768 -74
rect 1820 -126 1842 -74
rect 1894 -126 1900 -74
rect 1428 -127 1900 -126
tri 1530 -219 1622 -127 ne
rect 1622 -219 1900 -127
tri 1622 -251 1654 -219 ne
rect 1654 -378 1900 -219
tri 2308 -293 2382 -219 se
rect 2382 -241 2434 2005
tri 2382 -293 2434 -241 nw
tri 2234 -367 2308 -293 se
tri 2308 -367 2382 -293 nw
rect 2587 -297 2639 2436
tri 2639 2422 2653 2436 nw
rect 4046 733 4349 2684
tri 4848 2254 4958 2364 se
rect 4958 2332 5036 4354
tri 5036 4351 5039 4354 nw
tri 5816 4351 5819 4354 ne
rect 5819 4351 5906 4354
tri 5819 4316 5854 4351 ne
tri 5780 4021 5854 4095 se
rect 5854 4073 5906 4351
tri 5906 4316 5944 4354 nw
tri 5854 4021 5906 4073 nw
tri 5706 3947 5780 4021 se
tri 5780 3947 5854 4021 nw
tri 5667 3908 5706 3947 se
rect 5706 3908 5741 3947
tri 5741 3908 5780 3947 nw
tri 5632 3873 5667 3908 se
rect 5667 3873 5706 3908
tri 5706 3873 5741 3908 nw
tri 5615 3856 5632 3873 se
rect 5632 3856 5689 3873
tri 5689 3856 5706 3873 nw
tri 5558 3799 5615 3856 se
rect 5615 3799 5632 3856
tri 5632 3799 5689 3856 nw
tri 5484 3725 5558 3799 se
tri 5558 3725 5632 3799 nw
tri 5410 3651 5484 3725 se
tri 5484 3651 5558 3725 nw
tri 4958 2254 5036 2332 nw
tri 5397 3638 5410 3651 se
rect 5410 3638 5471 3651
tri 5471 3638 5484 3651 nw
tri 4738 2144 4848 2254 se
tri 4848 2144 4958 2254 nw
rect 4046 681 4052 733
rect 4104 681 4132 733
rect 4184 681 4212 733
rect 4264 681 4291 733
rect 4343 681 4349 733
rect 4046 659 4349 681
rect 4046 607 4052 659
rect 4104 607 4132 659
rect 4184 607 4212 659
rect 4264 607 4291 659
rect 4343 607 4349 659
rect 4046 585 4349 607
rect 4046 533 4052 585
rect 4104 533 4132 585
rect 4184 533 4212 585
rect 4264 533 4291 585
rect 4343 533 4349 585
rect 4046 20 4349 533
rect 4046 -32 4052 20
rect 4104 -32 4132 20
rect 4184 -32 4212 20
rect 4264 -32 4291 20
rect 4343 -32 4349 20
rect 4046 -74 4349 -32
rect 4046 -126 4052 -74
rect 4104 -126 4132 -74
rect 4184 -126 4212 -74
rect 4264 -126 4291 -74
rect 4343 -126 4349 -74
tri 2639 -297 2728 -208 sw
rect 2587 -318 2728 -297
tri 2728 -318 2749 -297 sw
rect 2587 -327 3611 -318
tri 2223 -378 2234 -367 se
rect 2234 -378 2297 -367
tri 2297 -378 2308 -367 nw
rect 1654 -430 1660 -378
rect 1712 -430 1751 -378
rect 1803 -430 1842 -378
rect 1894 -430 1900 -378
tri 2171 -430 2223 -378 se
rect 2223 -430 2245 -378
tri 2245 -430 2297 -378 nw
rect 2587 -383 3555 -327
rect 2587 -407 3611 -383
tri 2160 -441 2171 -430 se
rect 2171 -441 2234 -430
tri 2234 -441 2245 -430 nw
tri 2157 -444 2160 -441 se
rect 2160 -444 2231 -441
tri 2231 -444 2234 -441 nw
rect 2157 -463 2212 -444
tri 2212 -463 2231 -444 nw
rect 2587 -463 3555 -407
rect 4046 -378 4349 -126
tri 4700 2106 4738 2144 se
rect 4738 2106 4810 2144
tri 4810 2106 4848 2144 nw
rect 4700 -297 4778 2106
tri 4778 2074 4810 2106 nw
rect 5397 1385 5449 3638
tri 5449 3616 5471 3638 nw
rect 5768 3521 5774 3573
rect 5826 3521 5838 3573
rect 5890 3521 5896 3573
rect 5768 1963 5820 3521
tri 5820 3487 5854 3521 nw
rect 6258 2083 6310 6021
rect 7388 6032 7394 6084
rect 7446 6032 7458 6084
rect 7510 6032 7516 6084
tri 14220 6041 14263 6084 se
rect 14263 6075 14312 6084
rect 14263 6041 14278 6075
tri 14278 6041 14312 6075 nw
tri 14354 6580 14357 6583 se
rect 14357 6580 14408 6583
tri 14408 6580 14436 6608 nw
tri 14219 6040 14220 6041 se
rect 14220 6040 14277 6041
tri 14277 6040 14278 6041 nw
tri 14214 6035 14219 6040 se
rect 14219 6035 14272 6040
tri 14272 6035 14277 6040 nw
tri 14349 6035 14354 6040 se
rect 14354 6035 14392 6580
tri 14392 6564 14408 6580 nw
tri 14617 6242 14651 6276 se
rect 14651 6242 14688 15478
rect 14560 6190 14566 6242
rect 14618 6190 14630 6242
rect 14682 6190 14688 6242
tri 14722 6244 14728 6250 se
rect 14728 6244 14768 15511
rect 15128 15225 15168 15417
tri 14768 6244 14774 6250 sw
rect 14722 6238 14774 6244
rect 14722 6174 14774 6186
rect 14722 6116 14774 6122
tri 14802 6163 14808 6169 se
rect 14808 6163 14848 15225
tri 14848 6163 14854 6169 sw
rect 14802 6157 14854 6163
rect 14802 6093 14854 6105
tri 14886 6080 14888 6082 se
rect 14888 6080 14928 15225
tri 14928 6080 14930 6082 sw
rect 14802 6035 14854 6041
rect 14882 6074 14934 6080
tri 14211 6032 14214 6035 se
rect 14214 6032 14269 6035
tri 14269 6032 14272 6035 nw
tri 14346 6032 14349 6035 se
rect 14349 6032 14392 6035
rect 7388 6022 7464 6032
tri 7464 6022 7474 6032 nw
tri 14201 6022 14211 6032 se
rect 14211 6022 14259 6032
tri 14259 6022 14269 6032 nw
tri 14336 6022 14346 6032 se
rect 14346 6022 14392 6032
rect 7388 6016 7458 6022
tri 7458 6016 7464 6022 nw
tri 14195 6016 14201 6022 se
rect 14201 6016 14253 6022
tri 14253 6016 14259 6022 nw
tri 14330 6016 14336 6022 se
rect 14336 6020 14392 6022
rect 14336 6016 14382 6020
tri 7359 3578 7388 3607 se
rect 7388 3578 7440 6016
tri 7440 5998 7458 6016 nw
rect 8166 5964 8172 6016
rect 8224 5964 8236 6016
rect 8288 5964 8294 6016
tri 14189 6010 14195 6016 se
rect 14195 6010 14247 6016
tri 14247 6010 14253 6016 nw
tri 14324 6010 14330 6016 se
rect 14330 6010 14382 6016
tri 14382 6010 14392 6020 nw
rect 14882 6010 14934 6022
tri 14161 5982 14189 6010 se
rect 14189 5982 14219 6010
tri 14219 5982 14247 6010 nw
tri 14296 5982 14324 6010 se
rect 14324 5982 14354 6010
tri 14354 5982 14382 6010 nw
tri 14156 5977 14161 5982 se
rect 14161 5977 14214 5982
tri 14214 5977 14219 5982 nw
tri 14291 5977 14296 5982 se
rect 14296 5977 14330 5982
tri 14155 5976 14156 5977 se
rect 14156 5976 14213 5977
tri 14213 5976 14214 5977 nw
tri 14290 5976 14291 5977 se
rect 14291 5976 14330 5977
tri 12072 5964 12084 5976 se
rect 12084 5964 14201 5976
tri 14201 5964 14213 5976 nw
tri 14278 5964 14290 5976 se
rect 14290 5964 14330 5976
rect 8166 5958 8246 5964
tri 8246 5958 8252 5964 nw
tri 12066 5958 12072 5964 se
rect 12072 5958 14195 5964
tri 14195 5958 14201 5964 nw
tri 14272 5958 14278 5964 se
rect 14278 5958 14330 5964
tri 14330 5958 14354 5982 nw
rect 8166 5952 8240 5958
tri 8240 5952 8246 5958 nw
tri 12060 5952 12066 5958 se
rect 12066 5952 14189 5958
tri 14189 5952 14195 5958 nw
tri 14266 5952 14272 5958 se
rect 14272 5952 14324 5958
tri 14324 5952 14330 5958 nw
rect 14882 5952 14934 5958
tri 14962 6000 14968 6006 se
rect 14968 6000 15008 15225
tri 15008 6000 15014 6006 sw
rect 14962 5994 15014 6000
rect 8166 5942 8230 5952
tri 8230 5942 8240 5952 nw
tri 12050 5942 12060 5952 se
rect 12060 5942 14179 5952
tri 14179 5942 14189 5952 nw
tri 14256 5942 14266 5952 se
rect 14266 5942 14314 5952
tri 14314 5942 14324 5952 nw
rect 8166 5936 8224 5942
tri 8224 5936 8230 5942 nw
tri 12044 5936 12050 5942 se
rect 12050 5936 14173 5942
tri 14173 5936 14179 5942 nw
tri 14250 5936 14256 5942 se
rect 14256 5936 14302 5942
rect 7961 5722 7967 5774
rect 8019 5722 8031 5774
rect 8083 5722 8089 5774
tri 8020 5693 8049 5722 ne
rect 7635 4569 7641 4621
rect 7693 4569 7705 4621
rect 7757 4569 7763 4621
tri 7635 4563 7641 4569 ne
rect 7641 4563 7757 4569
tri 7757 4563 7763 4569 nw
tri 7641 4532 7672 4563 ne
rect 7672 4532 7726 4563
tri 7726 4532 7757 4563 nw
tri 7598 3697 7672 3771 se
rect 7672 3749 7724 4532
tri 7724 4530 7726 4532 nw
tri 7672 3697 7724 3749 nw
tri 7537 3636 7598 3697 se
rect 7598 3636 7665 3697
tri 7665 3690 7672 3697 nw
tri 7440 3578 7469 3607 sw
rect 7537 3578 7665 3636
tri 7354 3573 7359 3578 se
rect 7359 3573 7469 3578
tri 7469 3573 7474 3578 sw
rect 7350 3521 7356 3573
rect 7408 3521 7420 3573
rect 7472 3521 7478 3573
rect 7537 3526 7543 3578
rect 7595 3526 7607 3578
rect 7659 3526 7665 3578
tri 8047 3526 8049 3528 se
rect 8049 3526 8089 5722
tri 8042 3521 8047 3526 se
rect 8047 3521 8089 3526
tri 7975 3454 8042 3521 se
rect 8042 3494 8089 3521
rect 8042 3454 8049 3494
tri 8049 3454 8089 3494 nw
tri 7927 3406 7975 3454 se
rect 7975 3406 8001 3454
tri 8001 3406 8049 3454 nw
tri 7901 3380 7927 3406 se
rect 7927 3380 7975 3406
tri 7975 3380 8001 3406 nw
tri 7875 3354 7901 3380 se
rect 7901 3354 7949 3380
tri 7949 3354 7975 3380 nw
tri 7842 3321 7875 3354 se
rect 7875 3321 7916 3354
tri 7916 3321 7949 3354 nw
tri 7779 2220 7842 2283 se
rect 7842 2261 7894 3321
tri 7894 3299 7916 3321 nw
tri 8092 2346 8166 2420 se
rect 8166 2398 8218 5936
tri 8218 5930 8224 5936 nw
rect 9186 5884 9192 5936
rect 9244 5884 9256 5936
rect 9308 5884 9314 5936
tri 12038 5930 12044 5936 se
rect 12044 5930 12096 5936
tri 12096 5930 12102 5936 nw
tri 14244 5930 14250 5936 se
rect 14250 5930 14302 5936
tri 14302 5930 14314 5942 nw
rect 14962 5930 15014 5942
tri 12032 5924 12038 5930 se
rect 12038 5924 12090 5930
tri 12090 5924 12096 5930 nw
tri 14238 5924 14244 5930 se
rect 14244 5924 14296 5930
tri 14296 5924 14302 5930 nw
tri 12026 5918 12032 5924 se
rect 12032 5918 12084 5924
tri 12084 5918 12090 5924 nw
tri 14232 5918 14238 5924 se
rect 14238 5918 14270 5924
tri 12006 5898 12026 5918 se
rect 12026 5898 12064 5918
tri 12064 5898 12084 5918 nw
tri 14212 5898 14232 5918 se
rect 14232 5898 14270 5918
tri 14270 5898 14296 5924 nw
tri 11992 5884 12006 5898 se
rect 12006 5884 12050 5898
tri 12050 5884 12064 5898 nw
tri 12136 5884 12150 5898 se
rect 12150 5884 14250 5898
tri 9193 5878 9199 5884 ne
rect 9199 5878 9295 5884
tri 9295 5878 9301 5884 nw
tri 11986 5878 11992 5884 se
rect 11992 5878 12044 5884
tri 12044 5878 12050 5884 nw
tri 12130 5878 12136 5884 se
rect 12136 5878 14250 5884
tri 14250 5878 14270 5898 nw
tri 9199 5863 9214 5878 ne
rect 9214 5872 9289 5878
tri 9289 5872 9295 5878 nw
tri 11980 5872 11986 5878 se
rect 11986 5872 12038 5878
tri 12038 5872 12044 5878 nw
tri 12124 5872 12130 5878 se
rect 12130 5872 14244 5878
tri 14244 5872 14250 5878 nw
rect 14962 5872 15014 5878
tri 15042 5914 15048 5920 se
rect 15048 5914 15088 15225
tri 15088 5914 15094 5920 sw
rect 15042 5908 15094 5914
rect 9214 5863 9280 5872
tri 9280 5863 9289 5872 nw
tri 11972 5864 11980 5872 se
rect 11980 5864 12030 5872
tri 12030 5864 12038 5872 nw
tri 12123 5871 12124 5872 se
rect 12124 5871 14243 5872
tri 14243 5871 14244 5872 nw
rect 11972 5863 12029 5864
tri 12029 5863 12030 5864 nw
rect 12123 5863 14235 5871
tri 14235 5863 14243 5871 nw
tri 9214 5850 9227 5863 ne
tri 9193 3952 9227 3986 se
rect 9227 3952 9267 5863
tri 9267 5850 9280 5863 nw
rect 9967 5811 9973 5863
rect 10025 5811 10037 5863
rect 10089 5811 10095 5863
tri 11971 5811 11972 5812 se
rect 11972 5811 12024 5863
tri 12024 5858 12029 5863 nw
rect 12123 5858 14230 5863
tri 14230 5858 14235 5863 nw
rect 12123 5856 12288 5858
tri 12288 5856 12290 5858 nw
rect 12123 5844 12276 5856
tri 12276 5844 12288 5856 nw
rect 15042 5844 15094 5856
rect 12123 5830 12262 5844
tri 12262 5830 12276 5844 nw
tri 12024 5811 12025 5812 sw
tri 9967 5781 9997 5811 ne
tri 9155 3914 9193 3952 se
rect 9193 3914 9229 3952
tri 9229 3914 9267 3952 nw
tri 9149 3908 9155 3914 se
rect 9155 3908 9223 3914
tri 9223 3908 9229 3914 nw
tri 9097 3856 9149 3908 se
rect 9149 3856 9171 3908
tri 9171 3856 9223 3908 nw
tri 9081 3840 9097 3856 se
rect 9097 3840 9155 3856
tri 9155 3840 9171 3856 nw
tri 9007 3766 9081 3840 se
tri 9081 3766 9155 3840 nw
tri 8933 3692 9007 3766 se
tri 9007 3692 9081 3766 nw
tri 8859 3618 8933 3692 se
tri 8933 3618 9007 3692 nw
tri 8848 3607 8859 3618 se
rect 8859 3607 8922 3618
tri 8922 3607 8933 3618 nw
tri 8819 3578 8848 3607 se
rect 8848 3578 8893 3607
tri 8893 3578 8922 3607 nw
tri 8814 3573 8819 3578 se
rect 8819 3573 8888 3578
tri 8888 3573 8893 3578 nw
tri 8785 3544 8814 3573 se
rect 8814 3544 8859 3573
tri 8859 3544 8888 3573 nw
tri 8767 3526 8785 3544 se
rect 8785 3526 8841 3544
tri 8841 3526 8859 3544 nw
tri 8762 3521 8767 3526 se
rect 8767 3521 8836 3526
tri 8836 3521 8841 3526 nw
tri 8166 2346 8218 2398 nw
tri 8733 3492 8762 3521 se
rect 8762 3492 8785 3521
rect 7842 2220 7853 2261
tri 7853 2220 7894 2261 nw
tri 8032 2286 8092 2346 se
rect 8092 2286 8106 2346
tri 8106 2286 8166 2346 nw
rect 7779 1506 7831 2220
tri 7831 2198 7853 2220 nw
rect 8032 1972 8084 2286
tri 8084 2264 8106 2286 nw
rect 8733 1992 8785 3492
tri 8785 3470 8836 3521 nw
rect 9997 3406 10037 5811
tri 10037 5781 10067 5811 nw
tri 11941 5781 11971 5811 se
rect 11971 5781 12025 5811
tri 11938 5778 11941 5781 se
rect 11941 5778 12025 5781
tri 12025 5778 12058 5811 sw
rect 12123 5778 12129 5830
rect 12181 5778 12193 5830
rect 12245 5778 12251 5830
tri 12251 5819 12262 5830 nw
rect 12304 5778 12310 5830
rect 12362 5778 12374 5830
rect 12426 5778 12432 5830
rect 15042 5786 15094 5792
tri 11934 5774 11938 5778 se
rect 11938 5774 12058 5778
tri 12058 5774 12062 5778 sw
tri 12129 5774 12133 5778 ne
rect 12133 5774 12247 5778
tri 12247 5774 12251 5778 nw
tri 12310 5774 12314 5778 ne
rect 12314 5774 12402 5778
rect 11934 5722 11940 5774
rect 11992 5722 12004 5774
rect 12056 5722 12062 5774
tri 12133 5744 12163 5774 ne
tri 12131 5189 12163 5221 se
rect 12163 5197 12221 5774
tri 12221 5748 12247 5774 nw
tri 12314 5748 12340 5774 ne
rect 12340 5748 12402 5774
tri 12402 5748 12432 5778 nw
tri 12340 5744 12344 5748 ne
rect 12163 5189 12213 5197
tri 12213 5189 12221 5197 nw
tri 12262 5189 12344 5271 se
rect 12344 5247 12402 5748
tri 13687 5493 13698 5504 se
rect 13698 5493 14338 5504
tri 14338 5493 14349 5504 sw
tri 13624 5430 13687 5493 se
rect 13687 5452 14349 5493
rect 13687 5430 13698 5452
tri 13698 5430 13720 5452 nw
tri 14316 5430 14338 5452 ne
rect 14338 5430 14349 5452
tri 13613 5419 13624 5430 se
rect 13624 5419 13687 5430
tri 13687 5419 13698 5430 nw
tri 14338 5419 14349 5430 ne
tri 14349 5419 14423 5493 sw
tri 13550 5356 13613 5419 se
rect 13613 5356 13624 5419
tri 13624 5356 13687 5419 nw
tri 14349 5397 14371 5419 ne
tri 12344 5189 12402 5247 nw
tri 13503 5309 13550 5356 se
rect 13550 5309 13577 5356
tri 13577 5309 13624 5356 nw
tri 12081 5139 12131 5189 se
rect 12131 5148 12172 5189
tri 12172 5148 12213 5189 nw
tri 12221 5148 12262 5189 se
rect 12131 5139 12163 5148
tri 12163 5139 12172 5148 nw
tri 12212 5139 12221 5148 se
rect 12221 5139 12262 5148
tri 12049 5107 12081 5139 se
rect 12081 5107 12131 5139
tri 12131 5107 12163 5139 nw
tri 12180 5107 12212 5139 se
rect 12212 5107 12262 5139
tri 12262 5107 12344 5189 nw
tri 11999 5057 12049 5107 se
rect 12049 5090 12114 5107
tri 12114 5090 12131 5107 nw
tri 12163 5090 12180 5107 se
rect 12049 5057 12081 5090
tri 12081 5057 12114 5090 nw
tri 12130 5057 12163 5090 se
rect 12163 5057 12180 5090
tri 11967 5025 11999 5057 se
rect 11999 5025 12049 5057
tri 12049 5025 12081 5057 nw
tri 12098 5025 12130 5057 se
rect 12130 5025 12180 5057
tri 12180 5025 12262 5107 nw
tri 11917 4975 11967 5025 se
rect 11967 5008 12032 5025
tri 12032 5008 12049 5025 nw
tri 12081 5008 12098 5025 se
rect 11967 4975 11999 5008
tri 11999 4975 12032 5008 nw
tri 12048 4975 12081 5008 se
rect 12081 4975 12098 5008
tri 11885 4943 11917 4975 se
rect 11917 4943 11967 4975
tri 11967 4943 11999 4975 nw
tri 12016 4943 12048 4975 se
rect 12048 4943 12098 4975
tri 12098 4943 12180 5025 nw
tri 11835 4893 11885 4943 se
rect 11885 4926 11950 4943
tri 11950 4926 11967 4943 nw
tri 11999 4926 12016 4943 se
rect 11885 4893 11917 4926
tri 11917 4893 11950 4926 nw
tri 11966 4893 11999 4926 se
rect 11999 4893 12016 4926
tri 11803 4861 11835 4893 se
rect 11835 4861 11885 4893
tri 11885 4861 11917 4893 nw
tri 11934 4861 11966 4893 se
rect 11966 4861 12016 4893
tri 12016 4861 12098 4943 nw
tri 11753 4811 11803 4861 se
rect 11803 4844 11868 4861
tri 11868 4844 11885 4861 nw
tri 11917 4844 11934 4861 se
rect 11934 4844 11945 4861
rect 11803 4811 11835 4844
tri 11835 4811 11868 4844 nw
tri 11884 4811 11917 4844 se
rect 11917 4811 11945 4844
tri 11682 4740 11753 4811 se
rect 11753 4740 11764 4811
tri 11764 4740 11835 4811 nw
tri 11863 4790 11884 4811 se
rect 11884 4790 11945 4811
tri 11945 4790 12016 4861 nw
tri 11613 3908 11682 3977 se
rect 11682 3908 11741 4740
tri 11741 4717 11764 4740 nw
rect 10259 3856 10265 3908
rect 10317 3856 10329 3908
rect 10381 3856 10387 3908
rect 11613 3856 11619 3908
rect 11671 3856 11683 3908
rect 11735 3856 11741 3908
tri 10037 3406 10125 3494 sw
rect 9997 3354 10003 3406
rect 10055 3354 10067 3406
rect 10119 3354 10125 3406
tri 8733 1981 8744 1992 ne
rect 8744 1981 8785 1992
tri 8084 1972 8093 1981 sw
tri 8744 1972 8753 1981 ne
rect 8753 1972 8785 1981
tri 8785 1972 8827 2014 sw
rect 8032 1949 8093 1972
tri 8093 1949 8116 1972 sw
tri 8753 1949 8776 1972 ne
rect 8776 1949 8827 1972
tri 8827 1949 8850 1972 sw
rect 8032 1940 8116 1949
tri 8116 1940 8125 1949 sw
tri 8776 1940 8785 1949 ne
rect 8785 1940 8850 1949
rect 8032 1929 8125 1940
tri 8125 1929 8136 1940 sw
rect 8032 1878 8136 1929
tri 8785 1920 8805 1940 ne
rect 8805 1920 8850 1940
tri 8850 1920 8879 1949 sw
tri 8805 1908 8817 1920 ne
rect 8817 1908 8879 1920
tri 8879 1908 8891 1920 sw
tri 8032 1875 8035 1878 ne
rect 8035 1875 8136 1878
tri 8817 1875 8850 1908 ne
rect 8850 1875 8891 1908
tri 8891 1875 8924 1908 sw
tri 8035 1856 8054 1875 ne
rect 8054 1856 8136 1875
tri 8850 1856 8869 1875 ne
rect 8869 1856 8924 1875
tri 8924 1856 8943 1875 sw
tri 8054 1855 8055 1856 ne
rect 8055 1855 8136 1856
tri 8869 1855 8870 1856 ne
rect 8870 1855 8943 1856
tri 8943 1855 8944 1856 sw
tri 8055 1826 8084 1855 ne
tri 7831 1506 7853 1528 sw
tri 7779 1505 7780 1506 ne
rect 7780 1505 7853 1506
tri 7853 1505 7854 1506 sw
tri 7780 1483 7802 1505 ne
rect 7802 1498 7854 1505
tri 7854 1498 7861 1505 sw
rect 7802 1483 7861 1498
tri 7802 1476 7809 1483 ne
tri 5449 1385 5471 1407 sw
tri 5397 1340 5442 1385 ne
rect 5442 1340 5471 1385
tri 5471 1340 5516 1385 sw
tri 5442 1311 5471 1340 ne
rect 5471 1311 5516 1340
tri 5516 1311 5545 1340 sw
tri 5471 1288 5494 1311 ne
rect 5494 1288 5545 1311
tri 5545 1288 5568 1311 sw
tri 5494 1237 5545 1288 ne
rect 5545 1286 5568 1288
tri 5568 1286 5570 1288 sw
rect 5545 1237 5570 1286
tri 5570 1237 5619 1286 sw
tri 5545 1215 5567 1237 ne
rect 5567 1234 5619 1237
tri 5619 1234 5622 1237 sw
rect 5567 1215 5622 1234
tri 5567 1212 5570 1215 ne
rect 5570 398 5622 1215
tri 7799 1205 7809 1215 se
rect 7809 1205 7861 1483
rect 7799 1193 7861 1205
rect 7799 1192 7860 1193
tri 7860 1192 7861 1193 nw
rect 7799 711 7851 1192
tri 7851 1183 7860 1192 nw
tri 7851 711 7873 733 sw
tri 7799 669 7841 711 ne
rect 7841 691 7873 711
tri 7873 691 7893 711 sw
tri 7838 454 7841 457 se
rect 7841 454 7893 691
tri 7818 434 7838 454 se
rect 7838 434 7893 454
tri 7808 424 7818 434 se
rect 7818 424 7893 434
rect 6069 355 6075 407
rect 6127 355 6139 407
rect 6191 372 6197 407
tri 6197 372 6220 395 sw
rect 7765 372 7771 424
rect 7823 372 7835 424
rect 7887 372 7893 424
rect 6191 362 6220 372
tri 6220 362 6230 372 sw
rect 6191 355 6230 362
tri 6230 355 6237 362 sw
tri 6170 348 6177 355 ne
rect 6177 348 6237 355
tri 6237 348 6244 355 sw
rect 5570 334 5622 346
tri 6177 329 6196 348 ne
rect 6196 344 6244 348
tri 6244 344 6248 348 sw
rect 5570 276 5622 282
rect 4046 -430 4052 -378
rect 4104 -430 4132 -378
rect 4184 -430 4212 -378
rect 4264 -430 4291 -378
rect 4343 -430 4349 -378
rect 6196 -318 6248 344
tri 8050 312 8084 346 se
rect 8084 312 8136 1855
tri 8870 1801 8924 1855 ne
rect 8924 1801 8944 1855
tri 8944 1801 8998 1855 sw
tri 8924 1727 8998 1801 ne
tri 8998 1727 9072 1801 sw
tri 8998 1653 9072 1727 ne
tri 9072 1653 9146 1727 sw
tri 9072 1579 9146 1653 ne
tri 9146 1579 9220 1653 sw
tri 9146 1505 9220 1579 ne
tri 9220 1505 9294 1579 sw
tri 9220 1483 9242 1505 ne
tri 8136 312 8170 346 sw
tri 9208 312 9242 346 se
rect 9242 312 9294 1505
tri 10254 1238 10259 1243 se
rect 10259 1238 10311 3856
tri 10311 3822 10345 3856 nw
rect 11603 3526 11609 3578
rect 11661 3526 11673 3578
rect 11725 3526 11731 3578
tri 11613 3521 11618 3526 ne
rect 11618 3521 11726 3526
tri 11726 3521 11731 3526 nw
tri 11618 3493 11646 3521 ne
tri 11153 2913 11205 2965 se
rect 11205 2913 11260 2965
rect 11312 2913 11324 2965
rect 11376 2913 11382 2965
tri 11117 2877 11153 2913 se
rect 11153 2877 11157 2913
rect 11117 2279 11157 2877
tri 11157 2859 11211 2913 nw
tri 11117 2265 11131 2279 ne
rect 11131 2265 11157 2279
tri 11157 2265 11189 2297 sw
tri 11131 2239 11157 2265 ne
rect 11157 2239 11189 2265
tri 11157 2207 11189 2239 ne
tri 11189 2207 11247 2265 sw
tri 11189 2149 11247 2207 ne
tri 11247 2149 11305 2207 sw
tri 11247 2091 11305 2149 ne
tri 11305 2091 11363 2149 sw
tri 11305 2033 11363 2091 ne
tri 11363 2033 11421 2091 sw
tri 11363 2015 11381 2033 ne
rect 10814 1972 10866 1978
rect 10814 1908 10866 1920
rect 10814 1850 10866 1856
rect 11149 1855 11155 1907
rect 11207 1855 11219 1907
rect 11271 1855 11277 1907
rect 11149 1675 11196 1855
tri 11196 1775 11276 1855 nw
tri 11196 1675 11200 1679 sw
rect 11149 1660 11200 1675
tri 11149 1609 11200 1660 ne
tri 11200 1609 11266 1675 sw
tri 11200 1590 11219 1609 ne
tri 10225 1209 10254 1238 se
rect 10254 1209 10311 1238
rect 10181 1157 10311 1209
rect 10181 1154 10264 1157
tri 10264 1154 10267 1157 nw
rect 10181 1140 10250 1154
tri 10250 1140 10264 1154 nw
rect 10181 1126 10236 1140
tri 10236 1126 10250 1140 nw
rect 10181 772 10233 1126
tri 10233 1123 10236 1126 nw
rect 11219 1025 11266 1609
rect 11381 1085 11421 2033
rect 11646 1290 11698 3521
tri 11698 3493 11726 3521 nw
rect 11863 1929 11922 4790
tri 11922 4767 11945 4790 nw
tri 13438 4639 13503 4704 se
rect 13503 4682 13555 5309
tri 13555 5287 13577 5309 nw
rect 13503 4639 13512 4682
tri 13512 4639 13555 4682 nw
tri 13432 4633 13438 4639 se
rect 13438 4633 13506 4639
tri 13506 4633 13512 4639 nw
rect 14371 4633 14423 5419
tri 13429 4630 13432 4633 se
rect 13432 4630 13503 4633
tri 13503 4630 13506 4633 nw
tri 13398 4599 13429 4630 se
rect 13429 4599 13472 4630
tri 13472 4599 13503 4630 nw
tri 12553 4581 12571 4599 se
rect 12571 4581 13454 4599
tri 13454 4581 13472 4599 nw
tri 12535 4563 12553 4581 se
rect 12553 4563 13436 4581
tri 13436 4563 13454 4581 nw
rect 14371 4563 14423 4581
tri 12497 4525 12535 4563 se
rect 12535 4547 13420 4563
tri 13420 4547 13436 4563 nw
rect 12535 4525 12571 4547
tri 12571 4525 12593 4547 nw
tri 12483 4511 12497 4525 se
rect 12497 4511 12557 4525
tri 12557 4511 12571 4525 nw
tri 12477 4505 12483 4511 se
rect 12483 4505 12551 4511
tri 12551 4505 12557 4511 nw
rect 14371 4505 14423 4511
tri 12465 4493 12477 4505 se
rect 12477 4493 12539 4505
tri 12539 4493 12551 4505 nw
tri 12442 3822 12465 3845 se
rect 12465 3823 12517 4493
tri 12517 4471 12539 4493 nw
rect 12465 3822 12511 3823
tri 12437 3817 12442 3822 se
rect 12442 3817 12511 3822
tri 12511 3817 12517 3823 nw
rect 12437 3035 12489 3817
tri 12489 3795 12511 3817 nw
rect 12437 2971 12489 2983
rect 12437 2913 12489 2919
rect 14640 2790 14917 2796
rect 14640 2738 14642 2790
rect 14694 2738 14716 2790
rect 14768 2738 14790 2790
rect 14842 2738 14864 2790
rect 14916 2738 14917 2790
rect 14640 2715 14917 2738
rect 14640 2663 14642 2715
rect 14694 2663 14716 2715
rect 14768 2663 14790 2715
rect 14842 2663 14864 2715
rect 14916 2663 14917 2715
rect 14640 2640 14917 2663
rect 14640 2588 14642 2640
rect 14694 2588 14716 2640
rect 14768 2588 14790 2640
rect 14842 2588 14864 2640
rect 14916 2588 14917 2640
rect 14640 2564 14917 2588
rect 14640 2512 14642 2564
rect 14694 2512 14716 2564
rect 14768 2512 14790 2564
rect 14842 2512 14864 2564
rect 14916 2512 14917 2564
rect 14640 2488 14917 2512
rect 14640 2436 14642 2488
rect 14694 2436 14716 2488
rect 14768 2436 14790 2488
rect 14842 2436 14864 2488
rect 14916 2436 14917 2488
tri 11922 1929 11945 1952 sw
tri 11863 1890 11902 1929 ne
rect 11902 1913 11945 1929
tri 11945 1913 11961 1929 sw
tri 11872 1340 11902 1370 se
rect 11902 1340 11961 1913
tri 11646 1288 11648 1290 ne
rect 11648 1288 11698 1290
tri 11698 1288 11722 1312 sw
rect 11833 1288 11839 1340
rect 11891 1288 11903 1340
rect 11955 1288 11961 1340
tri 11648 1250 11686 1288 ne
rect 11686 1250 11722 1288
tri 11722 1250 11760 1288 sw
tri 11686 1238 11698 1250 ne
rect 11698 1238 11760 1250
tri 11698 1192 11744 1238 ne
rect 11744 1192 11760 1238
tri 11760 1192 11818 1250 sw
rect 12572 1192 12624 1198
tri 11744 1176 11760 1192 ne
rect 11760 1176 11818 1192
tri 11818 1176 11834 1192 sw
tri 11760 1154 11782 1176 ne
tri 11381 1083 11383 1085 ne
rect 11383 1083 11421 1085
tri 11421 1083 11441 1103 sw
tri 11383 1074 11392 1083 ne
rect 11392 1074 11441 1083
tri 11441 1074 11450 1083 sw
tri 11392 1045 11421 1074 ne
rect 11421 1045 11450 1074
tri 11421 1026 11440 1045 ne
rect 11440 1026 11450 1045
tri 11266 1025 11267 1026 sw
tri 11440 1025 11441 1026 ne
rect 11441 1025 11450 1026
tri 11450 1025 11499 1074 sw
rect 11219 997 11267 1025
tri 11219 967 11249 997 ne
rect 11249 967 11267 997
tri 11267 967 11325 1025 sw
tri 11441 967 11499 1025 ne
tri 11499 967 11557 1025 sw
tri 11249 950 11266 967 ne
rect 11266 950 11325 967
tri 11266 894 11322 950 ne
rect 11322 949 11325 950
tri 11325 949 11343 967 sw
tri 11499 949 11517 967 ne
rect 11322 894 11343 949
tri 11343 894 11398 949 sw
rect 11151 842 11157 894
rect 11209 842 11221 894
rect 11273 842 11279 894
tri 11322 891 11325 894 ne
rect 11325 891 11398 894
tri 11398 891 11401 894 sw
tri 11325 888 11328 891 ne
rect 11328 888 11401 891
tri 11328 867 11349 888 ne
rect 11151 836 11273 842
tri 11273 836 11279 842 nw
rect 11151 824 11261 836
tri 11261 824 11273 836 nw
tri 10233 772 10251 790 sw
rect 10181 756 10251 772
tri 10251 756 10267 772 sw
rect 11151 757 11257 824
tri 11257 820 11261 824 nw
rect 11151 756 11256 757
tri 11256 756 11257 757 nw
rect 10181 704 10311 756
tri 10225 670 10259 704 ne
tri 10256 382 10259 385 se
rect 10259 382 10311 704
tri 10236 362 10256 382 se
rect 10256 362 10311 382
tri 10222 348 10236 362 se
rect 10236 348 10311 362
tri 9294 312 9327 345 sw
rect 8045 260 8051 312
rect 8103 260 8117 312
rect 8169 260 8175 312
rect 9203 260 9209 312
rect 9261 260 9275 312
rect 9327 260 9333 312
rect 10183 296 10189 348
rect 10241 296 10253 348
rect 10305 296 10311 348
tri 6248 -318 6264 -302 sw
rect 6196 -324 6264 -318
tri 6264 -324 6270 -318 sw
tri 6196 -398 6270 -324 ne
tri 6270 -398 6344 -324 sw
tri 6270 -430 6302 -398 ne
rect 6302 -430 6344 -398
tri 6302 -463 6335 -430 ne
rect 6335 -451 6344 -430
tri 6344 -451 6397 -398 sw
rect 6335 -463 6397 -451
tri 6397 -463 6409 -451 sw
rect 2157 -626 2209 -463
tri 2209 -466 2212 -463 nw
rect 2587 -472 3611 -463
tri 6335 -472 6344 -463 ne
rect 6344 -472 6409 -463
tri 6409 -472 6418 -463 sw
tri 6344 -515 6387 -472 ne
rect 6387 -503 6418 -472
tri 6418 -503 6449 -472 sw
rect 6387 -515 6449 -503
tri 6387 -525 6397 -515 ne
rect 6397 -626 6449 -515
rect 10438 -515 10444 -463
rect 10496 -515 10508 -463
rect 10560 -515 10566 -463
tri 10438 -534 10457 -515 ne
rect 10457 -534 10520 -515
tri 10520 -534 10539 -515 nw
rect 10457 -543 10511 -534
tri 10511 -543 10520 -534 nw
rect 10457 -630 10509 -543
tri 10509 -545 10511 -543 nw
rect 10551 -595 10557 -543
rect 10609 -595 10621 -543
rect 10673 -595 10679 -543
rect 10551 -631 10603 -595
tri 10603 -629 10637 -595 nw
rect 11151 -630 11203 756
tri 11203 703 11256 756 nw
tri 11318 703 11349 734 se
rect 11349 712 11401 888
tri 11275 660 11318 703 se
rect 11318 660 11349 703
tri 11349 660 11401 712 nw
tri 11263 648 11275 660 se
rect 11275 648 11337 660
tri 11337 648 11349 660 nw
tri 11245 630 11263 648 se
rect 11263 630 11319 648
tri 11319 630 11337 648 nw
rect 11245 -630 11297 630
tri 11297 608 11319 630 nw
tri 2891 -2202 2914 -2179 se
rect 2914 -2202 3209 -2179
rect 2891 -2235 3209 -2202
rect 3265 -2235 3289 -2179
rect 3345 -2235 3354 -2179
tri 2853 -2634 2891 -2596 se
rect 2891 -2634 2943 -2235
tri 2943 -2282 2990 -2235 nw
tri 2943 -2634 2981 -2596 sw
rect 2853 -2686 2859 -2634
rect 2911 -2686 2923 -2634
rect 2975 -2686 2981 -2634
tri 11487 -2679 11517 -2649 se
rect 11517 -2679 11557 967
rect 11782 -632 11834 1176
rect 12572 1126 12624 1140
rect 12572 888 12624 1074
rect 12572 824 12624 836
rect 12572 735 12624 772
rect 14640 648 14917 2436
rect 14640 596 14642 648
rect 14694 596 14716 648
rect 14768 596 14790 648
rect 14842 596 14864 648
rect 14916 596 14917 648
rect 14640 577 14917 596
rect 14640 525 14642 577
rect 14694 525 14716 577
rect 14768 525 14790 577
rect 14842 525 14864 577
rect 14916 525 14917 577
rect 14640 506 14917 525
rect 14640 454 14642 506
rect 14694 454 14716 506
rect 14768 454 14790 506
rect 14842 454 14864 506
rect 14916 454 14917 506
rect 14640 434 14917 454
rect 14640 382 14642 434
rect 14694 382 14716 434
rect 14768 382 14790 434
rect 14842 382 14864 434
rect 14916 382 14917 434
rect 14640 362 14917 382
rect 14640 310 14642 362
rect 14694 310 14716 362
rect 14768 310 14790 362
rect 14842 310 14864 362
rect 14916 310 14917 362
rect 14640 304 14917 310
rect 12683 -256 12709 -207
rect 13154 -315 13203 -252
tri 13131 -451 13152 -430 se
rect 13152 -451 13204 -316
tri 13130 -452 13131 -451 se
rect 13131 -452 13204 -451
tri 13119 -463 13130 -452 se
rect 13130 -463 13193 -452
tri 13193 -463 13204 -452 nw
rect 12325 -515 12331 -463
rect 12383 -515 12395 -463
rect 12447 -515 13141 -463
tri 13141 -515 13193 -463 nw
tri 13227 -515 13237 -505 se
rect 13237 -515 13289 -316
rect 13322 -328 13371 -275
rect 13514 -373 13549 -328
rect 13686 -376 13720 -327
rect 14160 -371 14204 -322
tri 13430 -451 13504 -377 se
rect 13504 -439 13556 -376
tri 13504 -451 13516 -439 nw
tri 13418 -463 13430 -451 se
tri 13366 -515 13418 -463 se
rect 13418 -515 13430 -463
tri 13217 -525 13227 -515 se
rect 13227 -525 13289 -515
tri 13356 -525 13366 -515 se
rect 13366 -525 13430 -515
tri 13430 -525 13504 -451 nw
tri 13215 -527 13217 -525 se
rect 13217 -527 13289 -525
tri 13199 -543 13215 -527 se
rect 13215 -543 13273 -527
tri 13273 -543 13289 -527 nw
tri 13338 -543 13356 -525 se
rect 12325 -595 12331 -543
rect 12383 -595 12395 -543
rect 12447 -592 13224 -543
tri 13224 -592 13273 -543 nw
tri 13289 -592 13338 -543 se
rect 13338 -592 13356 -543
rect 12447 -595 13221 -592
tri 13221 -595 13224 -592 nw
tri 13286 -595 13289 -592 se
rect 13289 -595 13356 -592
tri 13282 -599 13286 -595 se
rect 13286 -599 13356 -595
tri 13356 -599 13430 -525 nw
tri 13271 -610 13282 -599 se
rect 13282 -610 13314 -599
tri 11782 -641 11791 -632 ne
rect 11791 -641 11834 -632
tri 11834 -641 11865 -610 sw
tri 13240 -641 13271 -610 se
rect 13271 -641 13314 -610
tri 13314 -641 13356 -599 nw
tri 11791 -684 11834 -641 ne
rect 11834 -684 13271 -641
tri 13271 -684 13314 -641 nw
tri 11834 -693 11843 -684 ne
rect 11843 -693 13262 -684
tri 13262 -693 13271 -684 nw
tri 11480 -2686 11487 -2679 se
rect 11487 -2686 11557 -2679
tri 11557 -2686 11564 -2679 sw
tri 11464 -2702 11480 -2686 se
rect 11480 -2702 11564 -2686
rect 11464 -2714 11564 -2702
tri 11564 -2714 11592 -2686 sw
rect 11464 -2766 11470 -2714
rect 11522 -2766 11534 -2714
rect 11586 -2766 11592 -2714
<< via2 >>
rect 3381 28591 3437 28647
rect 3515 28591 3571 28647
rect 3381 28509 3437 28565
rect 3515 28509 3571 28565
rect 3381 28427 3437 28483
rect 3515 28427 3571 28483
rect 3381 28345 3437 28401
rect 3515 28345 3571 28401
rect 3381 28263 3437 28319
rect 3515 28263 3571 28319
rect 3381 28181 3437 28237
rect 3515 28181 3571 28237
rect 3381 28099 3437 28155
rect 3515 28099 3571 28155
rect 3381 28017 3437 28073
rect 3515 28017 3571 28073
rect 3381 27935 3437 27991
rect 3515 27935 3571 27991
rect 3381 27853 3437 27909
rect 3515 27853 3571 27909
rect 3381 27771 3437 27827
rect 3515 27771 3571 27827
rect 3381 27689 3437 27745
rect 3515 27689 3571 27745
rect 3381 27606 3437 27662
rect 3515 27606 3571 27662
rect 3381 27523 3437 27579
rect 3515 27523 3571 27579
rect 5668 23586 5724 23642
rect 5812 23586 5868 23642
rect 5668 23514 5724 23548
rect 5812 23514 5868 23548
rect 5668 23492 5681 23514
rect 5681 23492 5724 23514
rect 5812 23492 5862 23514
rect 5862 23492 5868 23514
rect 5668 23440 5724 23453
rect 5812 23440 5868 23453
rect 5668 23397 5681 23440
rect 5681 23397 5724 23440
rect 5812 23397 5862 23440
rect 5862 23397 5868 23440
rect 3555 -383 3611 -327
rect 3555 -463 3611 -407
rect 3209 -2235 3265 -2179
rect 3289 -2235 3345 -2179
<< metal3 >>
rect 3373 28647 3583 28656
rect 3373 28591 3381 28647
rect 3437 28591 3515 28647
rect 3571 28591 3583 28647
rect 3373 28565 3583 28591
rect 3373 28509 3381 28565
rect 3437 28509 3515 28565
rect 3571 28509 3583 28565
rect 3373 28483 3583 28509
rect 3373 28427 3381 28483
rect 3437 28427 3515 28483
rect 3571 28427 3583 28483
rect 3373 28401 3583 28427
rect 3373 28345 3381 28401
rect 3437 28345 3515 28401
rect 3571 28345 3583 28401
rect 3373 28319 3583 28345
rect 3373 28263 3381 28319
rect 3437 28263 3515 28319
rect 3571 28263 3583 28319
rect 3373 28237 3583 28263
rect 3373 28181 3381 28237
rect 3437 28181 3515 28237
rect 3571 28181 3583 28237
rect 3373 28155 3583 28181
rect 3373 28099 3381 28155
rect 3437 28099 3515 28155
rect 3571 28099 3583 28155
rect 3373 28073 3583 28099
rect 3373 28017 3381 28073
rect 3437 28017 3515 28073
rect 3571 28017 3583 28073
rect 3373 27991 3583 28017
rect 3373 27935 3381 27991
rect 3437 27935 3515 27991
rect 3571 27935 3583 27991
rect 3373 27909 3583 27935
rect 3373 27853 3381 27909
rect 3437 27853 3515 27909
rect 3571 27853 3583 27909
rect 3373 27827 3583 27853
rect 3373 27771 3381 27827
rect 3437 27771 3515 27827
rect 3571 27771 3583 27827
rect 3373 27745 3583 27771
rect 3373 27689 3381 27745
rect 3437 27689 3515 27745
rect 3571 27689 3583 27745
rect 3373 27662 3583 27689
rect 3373 27606 3381 27662
rect 3437 27606 3515 27662
rect 3571 27606 3583 27662
rect 3373 27579 3583 27606
rect 3373 27523 3381 27579
rect 3437 27523 3515 27579
rect 3571 27523 3583 27579
rect 3373 25532 3583 27523
tri 3373 25336 3569 25532 ne
rect 3569 25336 3583 25532
tri 3583 25336 3867 25620 sw
tri 3569 25322 3583 25336 ne
rect 3583 25322 3867 25336
tri 3583 25038 3867 25322 ne
tri 3867 25038 4165 25336 sw
tri 3867 24889 4016 25038 ne
rect 4016 24889 4581 25038
tri 4581 24889 4730 25038 sw
tri 4016 24828 4077 24889 ne
rect 4077 24828 4730 24889
tri 4493 24591 4730 24828 ne
tri 4730 24591 5028 24889 sw
tri 4730 24503 4818 24591 ne
rect 4818 23959 5028 24591
tri 4818 23949 4828 23959 ne
rect 4828 23949 5028 23959
tri 5028 23949 5126 24047 sw
tri 4828 23749 5028 23949 ne
rect 5028 23749 5126 23949
tri 5028 23651 5126 23749 ne
tri 5126 23651 5424 23949 sw
tri 5126 23642 5135 23651 ne
rect 5135 23642 5873 23651
tri 5135 23586 5191 23642 ne
rect 5191 23586 5668 23642
rect 5724 23586 5812 23642
rect 5868 23586 5873 23642
tri 5191 23548 5229 23586 ne
rect 5229 23548 5873 23586
tri 5229 23492 5285 23548 ne
rect 5285 23492 5668 23548
rect 5724 23492 5812 23548
rect 5868 23492 5873 23548
tri 5285 23453 5324 23492 ne
rect 5324 23453 5873 23492
tri 5324 23397 5380 23453 ne
rect 5380 23397 5668 23453
rect 5724 23397 5812 23453
rect 5868 23397 5873 23453
tri 5380 23388 5389 23397 ne
rect 5389 23388 5873 23397
rect 3550 -327 3616 -322
rect 3550 -383 3555 -327
rect 3611 -383 3616 -327
rect 3550 -407 3616 -383
rect 3550 -463 3555 -407
rect 3611 -463 3616 -407
rect 3550 -642 3616 -463
tri 3550 -653 3561 -642 ne
rect 3561 -653 3616 -642
tri 3616 -653 3655 -614 sw
tri 3561 -708 3616 -653 ne
rect 3616 -708 3655 -653
tri 3616 -747 3655 -708 ne
tri 3655 -747 3749 -653 sw
tri 3655 -841 3749 -747 ne
tri 3749 -841 3843 -747 sw
tri 3749 -869 3777 -841 ne
tri 3749 -1681 3777 -1653 se
rect 3777 -1681 3843 -841
tri 3660 -1770 3749 -1681 se
rect 3749 -1770 3754 -1681
tri 3754 -1770 3843 -1681 nw
tri 3566 -1864 3660 -1770 se
tri 3660 -1864 3754 -1770 nw
tri 3472 -1958 3566 -1864 se
tri 3566 -1958 3660 -1864 nw
tri 3378 -2052 3472 -1958 se
tri 3472 -2052 3566 -1958 nw
tri 3284 -2146 3378 -2052 se
tri 3378 -2146 3472 -2052 nw
tri 3256 -2174 3284 -2146 se
rect 3284 -2174 3350 -2146
tri 3350 -2174 3378 -2146 nw
rect 3204 -2179 3350 -2174
rect 3204 -2235 3209 -2179
rect 3265 -2235 3289 -2179
rect 3345 -2235 3350 -2179
rect 3204 -2240 3350 -2235
use sky130_fd_io__gpio_odrvrv2  sky130_fd_io__gpio_odrvrv2_0
timestamp 1633016201
transform 1 0 100 0 1 15231
box -973 -13613 15198 16619
use sky130_fd_io__gpiov2_octl_dat  sky130_fd_io__gpiov2_octl_dat_0
timestamp 1633016201
transform 1 0 -103 0 1 -770
box -670 -1593 15418 8041
<< labels >>
flabel metal3 s 9295 30051 9295 30051 0 FreeSans 440 0 0 0 VGND_IO
port 1 nsew
flabel metal3 s 6572 30165 6572 30165 0 FreeSans 440 0 0 0 VGND_IO
port 1 nsew
flabel metal3 s 4983 30110 4983 30110 0 FreeSans 440 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 14375 4533 14418 4577 3 FreeSans 520 180 0 0 HLD_I_H_N
port 2 nsew
flabel metal1 s 14721 5357 14764 5395 3 FreeSans 520 180 0 0 OD_H
port 3 nsew
flabel metal1 s 14934 4574 15008 4609 3 FreeSans 520 180 0 0 SLOW
port 4 nsew
flabel metal1 s 14971 4591 14971 4591 3 FreeSans 520 180 0 0 SLOW
port 4 nsew
flabel metal1 s 14971 4591 14971 4591 3 FreeSans 520 180 0 0 SLOW
port 4 nsew
flabel metal1 s 14594 372 14905 604 3 FreeSans 520 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 14594 2490 14905 2722 3 FreeSans 520 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 13148 4040 13459 4215 3 FreeSans 520 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 12885 3938 12926 4139 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 185 3938 225 4140 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 12999 4019 13039 4221 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 205 4039 205 4039 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 185 532 227 734 3 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 185 -126 222 20 3 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 848 2683 890 2885 3 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 12531 2683 12573 2885 7 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 12536 -126 12573 20 7 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 12531 532 12573 734 7 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 206 633 206 633 3 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 203 -53 203 -53 3 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 869 2784 869 2784 3 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 12554 -53 12554 -53 7 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 14737 -509 14904 -353 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 14737 3488 14904 3644 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 13072 5034 13239 5190 3 FreeSans 520 180 0 0 VGND
port 6 nsew
flabel metal1 s 14737 1648 14904 1804 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 14820 3566 14820 3566 3 FreeSans 520 0 0 0 VGND
port 6 nsew
flabel metal1 s 12433 4188 12600 4285 3 FreeSans 520 180 0 0 VGND
port 6 nsew
flabel metal1 s 277 5087 317 5289 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 12797 4169 12837 4298 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 422 4168 462 4298 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 12999 5017 13039 5219 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 297 5188 297 5188 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 442 4233 442 4233 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 855 1542 897 1672 3 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 1150 2158 1192 2288 3 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 367 3209 409 3411 3 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 8924 3209 8966 3411 7 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 12054 2158 12096 2288 7 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 857 1058 899 1260 3 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 876 1607 876 1607 3 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 1171 2223 1171 2223 3 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 388 3310 388 3310 3 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 12031 2158 12073 2288 7 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 12155 1542 12197 1672 7 FreeSans 300 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 14751 5639 14886 5756 3 FreeSans 520 180 0 0 VPWR
port 7 nsew
flabel metal1 s 5832 5732 5899 6080 3 FreeSans 520 0 0 0 VPWR_KA
port 8 nsew
flabel metal1 s 13410 23185 13465 23518 3 FreeSans 520 0 0 0 PAD
port 9 nsew
flabel metal1 s 14264 15319 14340 15371 3 FreeSans 520 0 0 0 TIE_HI_ESD
port 10 nsew
flabel metal1 s 11900 15967 11932 16025 3 FreeSans 520 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 551 16163 1720 16308 3 FreeSans 520 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 4219 15407 5388 15552 3 FreeSans 520 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 2627 23516 2680 23562 3 FreeSans 520 0 0 0 VGND_IO
port 1 nsew
flabel metal1 s 529 14138 567 14205 3 FreeSans 520 270 0 0 VSSIO_AMX
port 11 nsew
flabel metal2 s 13154 -315 13203 -252 3 FreeSans 520 90 0 0 DM_H[0]
port 12 nsew
flabel metal2 s 13322 -328 13371 -275 3 FreeSans 520 90 0 0 DM_H[1]
port 13 nsew
flabel metal2 s 12683 -256 12709 -207 3 FreeSans 520 90 0 0 DM_H[2]
port 14 nsew
flabel metal2 s 14160 -371 14204 -322 3 FreeSans 520 90 0 0 DM_H_N[0]
port 15 nsew
flabel metal2 s 13686 -376 13720 -327 3 FreeSans 520 90 0 0 DM_H_N[1]
port 16 nsew
flabel metal2 s 13514 -373 13549 -328 3 FreeSans 520 90 0 0 DM_H_N[2]
port 17 nsew
flabel metal2 s 4723 -292 4761 -259 3 FreeSans 520 90 0 0 HLD_I_OVR_H
port 18 nsew
flabel metal2 s 3251 6108 3297 6154 7 FreeSans 300 0 0 0 OE_N
port 19 nsew
flabel metal2 s 3274 6131 3274 6131 7 FreeSans 300 0 0 0 OE_N
port 19 nsew
flabel metal2 s 3724 6115 3776 6154 3 FreeSans 520 0 0 0 OUT
port 20 nsew
flabel metal2 s 11216 19247 12757 20340 3 FreeSans 520 0 0 0 PAD
port 9 nsew
flabel metal2 s 11216 26085 12757 27178 3 FreeSans 520 0 0 0 PAD
port 9 nsew
flabel metal2 s 15128 15225 15168 15417 3 FreeSans 520 90 0 0 TIE_LO_ESD
port 21 nsew
flabel metal2 s 13427 17780 14596 18850 3 FreeSans 520 0 0 0 VCC_IO
port 5 nsew
flabel metal2 s 4626 27838 7525 28365 3 FreeSans 520 0 0 0 VGND_IO
port 1 nsew
flabel locali s 410 16553 502 16599 3 FreeSans 520 0 0 0 VGND
port 6 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 5749062
string GDS_START 5682886
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016076
<< checkpaint >>
rect -1270 -1270 2440 2440
<< pwell >>
rect -10 1090 1176 1176
rect -10 76 76 1090
rect 523 817 544 866
rect 1090 76 1176 1090
rect -10 -10 1176 76
<< locali >>
rect 16 1116 1150 1150
rect 16 50 50 1116
rect 1116 50 1150 1116
rect 16 16 1150 50
<< metal1 >>
rect 0 1068 66 1164
rect 0 1016 7 1068
rect 59 1016 66 1068
rect 0 988 66 1016
rect 0 936 7 988
rect 59 936 66 988
rect 0 908 66 936
rect 0 856 7 908
rect 59 856 66 908
rect 0 828 66 856
rect 0 776 7 828
rect 59 776 66 828
rect 0 748 66 776
rect 0 696 7 748
rect 59 696 66 748
rect 0 668 66 696
rect 0 616 7 668
rect 59 616 66 668
rect 0 588 66 616
rect 0 536 7 588
rect 59 536 66 588
rect 0 508 66 536
rect 0 456 7 508
rect 59 456 66 508
rect 0 428 66 456
rect 0 376 7 428
rect 59 376 66 428
rect 0 348 66 376
rect 0 296 7 348
rect 59 296 66 348
rect 0 268 66 296
rect 0 216 7 268
rect 59 216 66 268
rect 0 188 66 216
rect 0 136 7 188
rect 59 136 66 188
rect 0 66 66 136
rect 94 1159 1164 1164
rect 94 1107 147 1159
rect 199 1107 227 1159
rect 279 1107 307 1159
rect 359 1107 387 1159
rect 439 1107 467 1159
rect 519 1107 547 1159
rect 599 1107 627 1159
rect 679 1107 707 1159
rect 759 1107 787 1159
rect 839 1107 867 1159
rect 919 1107 947 1159
rect 999 1107 1027 1159
rect 1079 1107 1164 1159
rect 94 1102 1164 1107
rect 94 94 122 1102
rect 150 66 178 1074
rect 206 94 234 1102
rect 262 66 290 1074
rect 318 94 346 1102
rect 374 66 402 1074
rect 430 94 458 1102
rect 486 66 514 1074
rect 542 94 570 1102
rect 598 66 626 1074
rect 654 94 682 1102
rect 710 66 738 1074
rect 766 94 794 1102
rect 822 66 850 1074
rect 878 94 906 1102
rect 934 66 962 1074
rect 990 94 1018 1102
rect 1102 1079 1164 1102
rect 1046 66 1074 1074
rect 1102 1027 1107 1079
rect 1159 1027 1164 1079
rect 1102 999 1164 1027
rect 1102 947 1107 999
rect 1159 947 1164 999
rect 1102 919 1164 947
rect 1102 867 1107 919
rect 1159 867 1164 919
rect 1102 839 1164 867
rect 1102 787 1107 839
rect 1159 787 1164 839
rect 1102 759 1164 787
rect 1102 707 1107 759
rect 1159 707 1164 759
rect 1102 679 1164 707
rect 1102 627 1107 679
rect 1159 627 1164 679
rect 1102 599 1164 627
rect 1102 547 1107 599
rect 1159 547 1164 599
rect 1102 519 1164 547
rect 1102 467 1107 519
rect 1159 467 1164 519
rect 1102 439 1164 467
rect 1102 387 1107 439
rect 1159 387 1164 439
rect 1102 359 1164 387
rect 1102 307 1107 359
rect 1159 307 1164 359
rect 1102 279 1164 307
rect 1102 227 1107 279
rect 1159 227 1164 279
rect 1102 199 1164 227
rect 1102 147 1107 199
rect 1159 147 1164 199
rect 1102 94 1164 147
rect 0 59 1164 66
rect 0 7 56 59
rect 108 7 136 59
rect 188 7 216 59
rect 268 7 296 59
rect 348 7 376 59
rect 428 7 456 59
rect 508 7 536 59
rect 588 7 616 59
rect 668 7 696 59
rect 748 7 776 59
rect 828 7 856 59
rect 908 7 936 59
rect 988 7 1016 59
rect 1068 7 1164 59
rect 0 0 1164 7
<< via1 >>
rect 7 1016 59 1068
rect 7 936 59 988
rect 7 856 59 908
rect 7 776 59 828
rect 7 696 59 748
rect 7 616 59 668
rect 7 536 59 588
rect 7 456 59 508
rect 7 376 59 428
rect 7 296 59 348
rect 7 216 59 268
rect 7 136 59 188
rect 147 1107 199 1159
rect 227 1107 279 1159
rect 307 1107 359 1159
rect 387 1107 439 1159
rect 467 1107 519 1159
rect 547 1107 599 1159
rect 627 1107 679 1159
rect 707 1107 759 1159
rect 787 1107 839 1159
rect 867 1107 919 1159
rect 947 1107 999 1159
rect 1027 1107 1079 1159
rect 1107 1027 1159 1079
rect 1107 947 1159 999
rect 1107 867 1159 919
rect 1107 787 1159 839
rect 1107 707 1159 759
rect 1107 627 1159 679
rect 1107 547 1159 599
rect 1107 467 1159 519
rect 1107 387 1159 439
rect 1107 307 1159 359
rect 1107 227 1159 279
rect 1107 147 1159 199
rect 56 7 108 59
rect 136 7 188 59
rect 216 7 268 59
rect 296 7 348 59
rect 376 7 428 59
rect 456 7 508 59
rect 536 7 588 59
rect 616 7 668 59
rect 696 7 748 59
rect 776 7 828 59
rect 856 7 908 59
rect 936 7 988 59
rect 1016 7 1068 59
<< metal2 >>
rect 66 1161 1164 1164
rect 66 1105 97 1161
rect 153 1159 223 1161
rect 279 1159 349 1161
rect 405 1159 475 1161
rect 531 1159 601 1161
rect 657 1159 727 1161
rect 783 1159 853 1161
rect 909 1159 979 1161
rect 1035 1159 1164 1161
rect 199 1107 223 1159
rect 279 1107 307 1159
rect 439 1107 467 1159
rect 531 1107 547 1159
rect 599 1107 601 1159
rect 679 1107 707 1159
rect 783 1107 787 1159
rect 839 1107 853 1159
rect 919 1107 947 1159
rect 1079 1107 1164 1159
rect 153 1105 223 1107
rect 279 1105 349 1107
rect 405 1105 475 1107
rect 531 1105 601 1107
rect 657 1105 727 1107
rect 783 1105 853 1107
rect 909 1105 979 1107
rect 1035 1105 1164 1107
rect 66 1102 1164 1105
rect 1102 1079 1164 1102
rect 0 1068 1074 1074
rect 0 1016 7 1068
rect 59 1046 1074 1068
rect 59 1016 66 1046
rect 1102 1035 1107 1079
rect 1159 1035 1164 1079
rect 1102 1018 1105 1035
rect 0 960 5 1016
rect 61 962 66 1016
rect 94 990 1105 1018
rect 1102 979 1105 990
rect 1161 979 1164 1035
rect 61 960 1074 962
rect 0 936 7 960
rect 59 936 1074 960
rect 0 934 1074 936
rect 1102 947 1107 979
rect 1159 947 1164 979
rect 0 908 66 934
rect 0 890 7 908
rect 59 890 66 908
rect 1102 919 1164 947
rect 1102 909 1107 919
rect 1159 909 1164 919
rect 1102 906 1105 909
rect 0 834 5 890
rect 61 850 66 890
rect 94 878 1105 906
rect 1102 853 1105 878
rect 1161 853 1164 909
rect 61 834 1074 850
rect 0 828 1074 834
rect 0 776 7 828
rect 59 822 1074 828
rect 1102 839 1164 853
rect 59 776 66 822
rect 1102 794 1107 839
rect 0 764 66 776
rect 94 787 1107 794
rect 1159 787 1164 839
rect 94 783 1164 787
rect 94 766 1105 783
rect 0 708 5 764
rect 61 738 66 764
rect 61 710 1074 738
rect 1102 727 1105 766
rect 1161 727 1164 783
rect 61 708 66 710
rect 0 696 7 708
rect 59 696 66 708
rect 0 668 66 696
rect 1102 707 1107 727
rect 1159 707 1164 727
rect 1102 682 1164 707
rect 0 638 7 668
rect 59 638 66 668
rect 94 679 1164 682
rect 94 657 1107 679
rect 1159 657 1164 679
rect 94 654 1105 657
rect 0 582 5 638
rect 61 626 66 638
rect 61 598 1074 626
rect 1102 601 1105 654
rect 1161 601 1164 657
rect 1102 599 1164 601
rect 61 582 66 598
rect 0 536 7 582
rect 59 536 66 582
rect 1102 570 1107 599
rect 94 547 1107 570
rect 1159 547 1164 599
rect 94 542 1164 547
rect 0 514 66 536
rect 1102 531 1164 542
rect 0 512 1074 514
rect 0 456 5 512
rect 61 486 1074 512
rect 61 456 66 486
rect 1102 475 1105 531
rect 1161 475 1164 531
rect 1102 467 1107 475
rect 1159 467 1164 475
rect 1102 458 1164 467
rect 0 428 66 456
rect 94 439 1164 458
rect 94 430 1107 439
rect 0 386 7 428
rect 59 402 66 428
rect 1102 405 1107 430
rect 1159 405 1164 439
rect 59 386 1074 402
rect 0 330 5 386
rect 61 374 1074 386
rect 61 330 66 374
rect 1102 349 1105 405
rect 1161 349 1164 405
rect 1102 346 1107 349
rect 0 296 7 330
rect 59 296 66 330
rect 94 318 1107 346
rect 0 290 66 296
rect 1102 307 1107 318
rect 1159 307 1164 349
rect 0 268 1074 290
rect 0 260 7 268
rect 59 262 1074 268
rect 1102 279 1164 307
rect 59 260 66 262
rect 0 204 5 260
rect 61 204 66 260
rect 1102 234 1105 279
rect 94 223 1105 234
rect 1161 223 1164 279
rect 94 206 1164 223
rect 0 188 66 204
rect 0 136 7 188
rect 59 178 66 188
rect 1102 199 1164 206
rect 59 150 1074 178
rect 1102 153 1107 199
rect 1159 153 1164 199
rect 59 136 66 150
rect 0 134 66 136
rect 0 78 5 134
rect 61 78 66 134
rect 1102 122 1105 153
rect 94 97 1105 122
rect 1161 97 1164 153
rect 94 94 1164 97
rect 0 66 66 78
rect 1102 66 1164 94
rect 0 61 1074 66
rect 0 59 78 61
rect 134 59 204 61
rect 260 59 330 61
rect 386 59 456 61
rect 512 59 582 61
rect 638 59 708 61
rect 764 59 834 61
rect 890 59 960 61
rect 1016 59 1074 61
rect 0 7 56 59
rect 134 7 136 59
rect 188 7 204 59
rect 268 7 296 59
rect 428 7 456 59
rect 512 7 536 59
rect 668 7 696 59
rect 764 7 776 59
rect 828 7 834 59
rect 908 7 936 59
rect 1068 7 1074 59
rect 0 5 78 7
rect 134 5 204 7
rect 260 5 330 7
rect 386 5 456 7
rect 512 5 582 7
rect 638 5 708 7
rect 764 5 834 7
rect 890 5 960 7
rect 1016 5 1074 7
rect 0 0 1074 5
<< via2 >>
rect 97 1159 153 1161
rect 223 1159 279 1161
rect 349 1159 405 1161
rect 475 1159 531 1161
rect 601 1159 657 1161
rect 727 1159 783 1161
rect 853 1159 909 1161
rect 979 1159 1035 1161
rect 97 1107 147 1159
rect 147 1107 153 1159
rect 223 1107 227 1159
rect 227 1107 279 1159
rect 349 1107 359 1159
rect 359 1107 387 1159
rect 387 1107 405 1159
rect 475 1107 519 1159
rect 519 1107 531 1159
rect 601 1107 627 1159
rect 627 1107 657 1159
rect 727 1107 759 1159
rect 759 1107 783 1159
rect 853 1107 867 1159
rect 867 1107 909 1159
rect 979 1107 999 1159
rect 999 1107 1027 1159
rect 1027 1107 1035 1159
rect 97 1105 153 1107
rect 223 1105 279 1107
rect 349 1105 405 1107
rect 475 1105 531 1107
rect 601 1105 657 1107
rect 727 1105 783 1107
rect 853 1105 909 1107
rect 979 1105 1035 1107
rect 1105 1027 1107 1035
rect 1107 1027 1159 1035
rect 1159 1027 1161 1035
rect 5 988 61 1016
rect 5 960 7 988
rect 7 960 59 988
rect 59 960 61 988
rect 1105 999 1161 1027
rect 1105 979 1107 999
rect 1107 979 1159 999
rect 1159 979 1161 999
rect 5 856 7 890
rect 7 856 59 890
rect 59 856 61 890
rect 5 834 61 856
rect 1105 867 1107 909
rect 1107 867 1159 909
rect 1159 867 1161 909
rect 1105 853 1161 867
rect 5 748 61 764
rect 5 708 7 748
rect 7 708 59 748
rect 59 708 61 748
rect 1105 759 1161 783
rect 1105 727 1107 759
rect 1107 727 1159 759
rect 1159 727 1161 759
rect 5 616 7 638
rect 7 616 59 638
rect 59 616 61 638
rect 5 588 61 616
rect 1105 627 1107 657
rect 1107 627 1159 657
rect 1159 627 1161 657
rect 1105 601 1161 627
rect 5 582 7 588
rect 7 582 59 588
rect 59 582 61 588
rect 5 508 61 512
rect 5 456 7 508
rect 7 456 59 508
rect 59 456 61 508
rect 1105 519 1161 531
rect 1105 475 1107 519
rect 1107 475 1159 519
rect 1159 475 1161 519
rect 5 376 7 386
rect 7 376 59 386
rect 59 376 61 386
rect 5 348 61 376
rect 5 330 7 348
rect 7 330 59 348
rect 59 330 61 348
rect 1105 387 1107 405
rect 1107 387 1159 405
rect 1159 387 1161 405
rect 1105 359 1161 387
rect 1105 349 1107 359
rect 1107 349 1159 359
rect 1159 349 1161 359
rect 5 216 7 260
rect 7 216 59 260
rect 59 216 61 260
rect 5 204 61 216
rect 1105 227 1107 279
rect 1107 227 1159 279
rect 1159 227 1161 279
rect 1105 223 1161 227
rect 5 78 61 134
rect 1105 147 1107 153
rect 1107 147 1159 153
rect 1159 147 1161 153
rect 1105 97 1161 147
rect 78 59 134 61
rect 204 59 260 61
rect 330 59 386 61
rect 456 59 512 61
rect 582 59 638 61
rect 708 59 764 61
rect 834 59 890 61
rect 960 59 1016 61
rect 78 7 108 59
rect 108 7 134 59
rect 204 7 216 59
rect 216 7 260 59
rect 330 7 348 59
rect 348 7 376 59
rect 376 7 386 59
rect 456 7 508 59
rect 508 7 512 59
rect 582 7 588 59
rect 588 7 616 59
rect 616 7 638 59
rect 708 7 748 59
rect 748 7 764 59
rect 834 7 856 59
rect 856 7 890 59
rect 960 7 988 59
rect 988 7 1016 59
rect 78 5 134 7
rect 204 5 260 7
rect 330 5 386 7
rect 456 5 512 7
rect 582 5 638 7
rect 708 5 764 7
rect 834 5 890 7
rect 960 5 1016 7
<< metal3 >>
rect 66 1165 1180 1180
rect 66 1161 219 1165
rect 66 1105 97 1161
rect 153 1105 219 1161
rect 66 1101 219 1105
rect 283 1101 345 1165
rect 409 1101 471 1165
rect 535 1101 597 1165
rect 661 1101 723 1165
rect 787 1101 849 1165
rect 913 1101 975 1165
rect 1039 1101 1101 1165
rect 1165 1101 1180 1165
rect 66 1086 1180 1101
rect 0 1020 66 1026
rect 0 956 1 1020
rect 65 956 66 1020
rect 0 894 66 956
rect 0 830 1 894
rect 65 830 66 894
rect 0 768 66 830
rect 0 704 1 768
rect 65 704 66 768
rect 0 642 66 704
rect 0 578 1 642
rect 65 578 66 642
rect 0 516 66 578
rect 0 452 1 516
rect 65 452 66 516
rect 0 390 66 452
rect 0 326 1 390
rect 65 326 66 390
rect 0 264 66 326
rect 0 200 1 264
rect 65 200 66 264
rect 0 138 66 200
rect 0 74 1 138
rect 65 74 66 138
rect 126 126 186 1086
rect 0 66 66 74
rect 246 66 306 1026
rect 366 126 426 1086
rect 486 66 546 1026
rect 606 126 666 1086
rect 726 66 786 1026
rect 846 126 906 1086
rect 1086 1039 1180 1086
rect 966 66 1026 1026
rect 1086 975 1101 1039
rect 1165 975 1180 1039
rect 1086 913 1180 975
rect 1086 849 1101 913
rect 1165 849 1180 913
rect 1086 787 1180 849
rect 1086 723 1101 787
rect 1165 723 1180 787
rect 1086 661 1180 723
rect 1086 597 1101 661
rect 1165 597 1180 661
rect 1086 535 1180 597
rect 1086 471 1101 535
rect 1165 471 1180 535
rect 1086 409 1180 471
rect 1086 345 1101 409
rect 1165 345 1180 409
rect 1086 283 1180 345
rect 1086 219 1101 283
rect 1165 219 1180 283
rect 1086 153 1180 219
rect 1086 97 1105 153
rect 1161 97 1180 153
rect 1086 66 1180 97
rect 0 65 1026 66
rect 0 1 74 65
rect 138 1 200 65
rect 264 1 326 65
rect 390 1 452 65
rect 516 1 578 65
rect 642 1 704 65
rect 768 1 830 65
rect 894 1 956 65
rect 1020 1 1026 65
rect 0 0 1026 1
<< via3 >>
rect 219 1161 283 1165
rect 219 1105 223 1161
rect 223 1105 279 1161
rect 279 1105 283 1161
rect 219 1101 283 1105
rect 345 1161 409 1165
rect 345 1105 349 1161
rect 349 1105 405 1161
rect 405 1105 409 1161
rect 345 1101 409 1105
rect 471 1161 535 1165
rect 471 1105 475 1161
rect 475 1105 531 1161
rect 531 1105 535 1161
rect 471 1101 535 1105
rect 597 1161 661 1165
rect 597 1105 601 1161
rect 601 1105 657 1161
rect 657 1105 661 1161
rect 597 1101 661 1105
rect 723 1161 787 1165
rect 723 1105 727 1161
rect 727 1105 783 1161
rect 783 1105 787 1161
rect 723 1101 787 1105
rect 849 1161 913 1165
rect 849 1105 853 1161
rect 853 1105 909 1161
rect 909 1105 913 1161
rect 849 1101 913 1105
rect 975 1161 1039 1165
rect 975 1105 979 1161
rect 979 1105 1035 1161
rect 1035 1105 1039 1161
rect 975 1101 1039 1105
rect 1101 1101 1165 1165
rect 1 1016 65 1020
rect 1 960 5 1016
rect 5 960 61 1016
rect 61 960 65 1016
rect 1 956 65 960
rect 1 890 65 894
rect 1 834 5 890
rect 5 834 61 890
rect 61 834 65 890
rect 1 830 65 834
rect 1 764 65 768
rect 1 708 5 764
rect 5 708 61 764
rect 61 708 65 764
rect 1 704 65 708
rect 1 638 65 642
rect 1 582 5 638
rect 5 582 61 638
rect 61 582 65 638
rect 1 578 65 582
rect 1 512 65 516
rect 1 456 5 512
rect 5 456 61 512
rect 61 456 65 512
rect 1 452 65 456
rect 1 386 65 390
rect 1 330 5 386
rect 5 330 61 386
rect 61 330 65 386
rect 1 326 65 330
rect 1 260 65 264
rect 1 204 5 260
rect 5 204 61 260
rect 61 204 65 260
rect 1 200 65 204
rect 1 134 65 138
rect 1 78 5 134
rect 5 78 61 134
rect 61 78 65 134
rect 1 74 65 78
rect 1101 1035 1165 1039
rect 1101 979 1105 1035
rect 1105 979 1161 1035
rect 1161 979 1165 1035
rect 1101 975 1165 979
rect 1101 909 1165 913
rect 1101 853 1105 909
rect 1105 853 1161 909
rect 1161 853 1165 909
rect 1101 849 1165 853
rect 1101 783 1165 787
rect 1101 727 1105 783
rect 1105 727 1161 783
rect 1161 727 1165 783
rect 1101 723 1165 727
rect 1101 657 1165 661
rect 1101 601 1105 657
rect 1105 601 1161 657
rect 1161 601 1165 657
rect 1101 597 1165 601
rect 1101 531 1165 535
rect 1101 475 1105 531
rect 1105 475 1161 531
rect 1161 475 1165 531
rect 1101 471 1165 475
rect 1101 405 1165 409
rect 1101 349 1105 405
rect 1105 349 1161 405
rect 1161 349 1165 405
rect 1101 345 1165 349
rect 1101 279 1165 283
rect 1101 223 1105 279
rect 1105 223 1161 279
rect 1161 223 1165 279
rect 1101 219 1165 223
rect 74 61 138 65
rect 74 5 78 61
rect 78 5 134 61
rect 134 5 138 61
rect 74 1 138 5
rect 200 61 264 65
rect 200 5 204 61
rect 204 5 260 61
rect 260 5 264 61
rect 200 1 264 5
rect 326 61 390 65
rect 326 5 330 61
rect 330 5 386 61
rect 386 5 390 61
rect 326 1 390 5
rect 452 61 516 65
rect 452 5 456 61
rect 456 5 512 61
rect 512 5 516 61
rect 452 1 516 5
rect 578 61 642 65
rect 578 5 582 61
rect 582 5 638 61
rect 638 5 642 61
rect 578 1 642 5
rect 704 61 768 65
rect 704 5 708 61
rect 708 5 764 61
rect 764 5 768 61
rect 704 1 768 5
rect 830 61 894 65
rect 830 5 834 61
rect 834 5 890 61
rect 890 5 894 61
rect 830 1 894 5
rect 956 61 1020 65
rect 956 5 960 61
rect 960 5 1016 61
rect 1016 5 1020 61
rect 956 1 1020 5
<< metal4 >>
rect 0 1026 66 1180
rect 126 1165 1180 1180
rect 126 1101 219 1165
rect 283 1101 345 1165
rect 409 1101 471 1165
rect 535 1101 597 1165
rect 661 1101 723 1165
rect 787 1101 849 1165
rect 913 1101 975 1165
rect 1039 1101 1101 1165
rect 1165 1101 1180 1165
rect 126 1086 1180 1101
rect 1086 1039 1180 1086
rect 0 1020 1026 1026
rect 0 956 1 1020
rect 65 966 1026 1020
rect 1086 975 1101 1039
rect 1165 975 1180 1039
rect 65 956 66 966
rect 0 894 66 956
rect 1086 913 1180 975
rect 1086 906 1101 913
rect 0 830 1 894
rect 65 830 66 894
rect 126 849 1101 906
rect 1165 849 1180 913
rect 126 846 1180 849
rect 0 786 66 830
rect 1086 787 1180 846
rect 0 768 1026 786
rect 0 704 1 768
rect 65 726 1026 768
rect 65 704 66 726
rect 0 642 66 704
rect 1086 723 1101 787
rect 1165 723 1180 787
rect 1086 666 1180 723
rect 0 578 1 642
rect 65 578 66 642
rect 126 661 1180 666
rect 126 606 1101 661
rect 0 546 66 578
rect 1086 597 1101 606
rect 1165 597 1180 661
rect 0 516 1026 546
rect 0 452 1 516
rect 65 486 1026 516
rect 1086 535 1180 597
rect 65 452 66 486
rect 0 390 66 452
rect 1086 471 1101 535
rect 1165 471 1180 535
rect 1086 426 1180 471
rect 0 326 1 390
rect 65 326 66 390
rect 126 409 1180 426
rect 126 366 1101 409
rect 0 306 66 326
rect 1086 345 1101 366
rect 1165 345 1180 409
rect 0 264 1026 306
rect 0 200 1 264
rect 65 246 1026 264
rect 1086 283 1180 345
rect 65 200 66 246
rect 0 138 66 200
rect 1086 219 1101 283
rect 1165 219 1180 283
rect 1086 186 1180 219
rect 0 74 1 138
rect 65 74 66 138
rect 126 126 1180 186
rect 0 66 66 74
rect 0 65 1180 66
rect 0 1 74 65
rect 138 1 200 65
rect 264 1 326 65
rect 390 1 452 65
rect 516 1 578 65
rect 642 1 704 65
rect 768 1 830 65
rect 894 1 956 65
rect 1020 1 1180 65
rect 0 0 1180 1
<< labels >>
flabel metal2 s 457 432 493 456 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel metal2 s 422 491 441 511 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel pwell s 523 817 544 866 0 FreeSans 400 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 202044
string GDS_START 187900
string path 28.750 28.325 0.400 28.325 
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1288 -1260 3416 1731
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_0
timestamp 1633016201
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_1
timestamp 1633016201
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_2
timestamp 1633016201
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_3
timestamp 1633016201
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_4
timestamp 1633016201
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_5
timestamp 1633016201
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_6
timestamp 1633016201
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_7
timestamp 1633016201
transform 1 0 1036 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_8
timestamp 1633016201
transform 1 0 1192 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_9
timestamp 1633016201
transform 1 0 1348 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_10
timestamp 1633016201
transform 1 0 1504 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_11
timestamp 1633016201
transform 1 0 1660 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_12
timestamp 1633016201
transform 1 0 1816 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_13
timestamp 1633016201
transform 1 0 1972 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_14
timestamp 1633016201
transform 1 0 2128 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 2156 471 2156 471 0 FreeSans 300 0 0 0 S
flabel comment s 2000 471 2000 471 0 FreeSans 300 0 0 0 D
flabel comment s 1844 471 1844 471 0 FreeSans 300 0 0 0 S
flabel comment s 1688 471 1688 471 0 FreeSans 300 0 0 0 D
flabel comment s 1532 471 1532 471 0 FreeSans 300 0 0 0 S
flabel comment s 1376 471 1376 471 0 FreeSans 300 0 0 0 D
flabel comment s 1220 471 1220 471 0 FreeSans 300 0 0 0 S
flabel comment s 1064 471 1064 471 0 FreeSans 300 0 0 0 D
flabel comment s 908 471 908 471 0 FreeSans 300 0 0 0 S
flabel comment s 752 471 752 471 0 FreeSans 300 0 0 0 D
flabel comment s 596 471 596 471 0 FreeSans 300 0 0 0 S
flabel comment s 440 471 440 471 0 FreeSans 300 0 0 0 D
flabel comment s 284 471 284 471 0 FreeSans 300 0 0 0 S
flabel comment s 128 471 128 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 27102
string GDS_START 19438
<< end >>

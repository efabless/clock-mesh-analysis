
VVDD      vpwr_0 0  1.8
VNB       VNB  0  0
VVGND     VGND 0  0

RP_clk_buf1_0 vpwr_0 vpwr_clk_buf1_branch_0  10
RP_clk_buf1_1 vpwr_0 vpwr_clk_buf1_branch_1  10
RP_clk_buf1_2 vpwr_0 vpwr_clk_buf1_branch_2  10
RP_clk_buf1_3 vpwr_0 vpwr_clk_buf1_branch_3  10
RP_clk_buf1_4 vpwr_0 vpwr_clk_buf1_branch_4  10
RP_clk_buf1_5 vpwr_0 vpwr_clk_buf1_branch_5  10
RP_clk_buf1_6 vpwr_0 vpwr_clk_buf1_branch_6  10
RP_clk_buf1_LOAD_0  vpwr_clk_buf1_branch_0 vpwr_clk_buf1_0 50
RP_clk_buf1_LOAD_1  vpwr_clk_buf1_branch_1 vpwr_clk_buf1_1 50
XDC_clk_buf1_0_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_3_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_4_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_5_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_6_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_7_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_8_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_9_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_10_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_11_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_12_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_13_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_14_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_15_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_16_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_17_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_18_0 VGND VNB vpwr_clk_buf1_0 vpwr_clk_buf1_0 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_0_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_1_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_2_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_3_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_4_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_5_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_6_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_7_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_8_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_9_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_10_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_11_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_12_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_13_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_14_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_15_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_16_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_17_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12
XDC_clk_buf1_18_1 VGND VNB vpwr_clk_buf1_1 vpwr_clk_buf1_1 sky130_fd_sc_hd__decap_12

VC_0  clk_0  VGND pulse 0 1.8 1.57n 1n 1n 48n 100n
VC_1  clk_1  VGND pulse 0 1.8 0.19n 1n 1n 48n 100n

x1_0  clk_0  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  co_0  sky130_fd_sc_hd__clkbuf_1
x1_1  clk_1  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  co_1  sky130_fd_sc_hd__clkbuf_1

R_0  co_0  co_1  70
R_1  co_1  co_2  70

x_buf1_buf16_intcon_0_0  co_0 co_i_0_0  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_1  co_0 co_i_0_1  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_2  co_0 co_i_0_2  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_3  co_0 co_i_0_3  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_4  co_0 co_i_0_4  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_5  co_0 co_i_0_5  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_6  co_0 co_i_0_6  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_7  co_0 co_i_0_7  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_8  co_0 co_i_0_8  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_9  co_0 co_i_0_9  VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_10 co_0 co_i_0_10 VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_11 co_0 co_i_0_11 VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_12 co_0 co_i_0_12 VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_13 co_0 co_i_0_13 VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_14 co_0 co_i_0_14 VGND int_con C=8f R=120
x_buf1_buf16_intcon_0_15 co_0 co_i_0_15 VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_0  co_1 co_i_1_0  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_1  co_1 co_i_1_1  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_2  co_1 co_i_1_2  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_3  co_1 co_i_1_3  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_4  co_1 co_i_1_4  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_5  co_1 co_i_1_5  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_6  co_1 co_i_1_6  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_7  co_1 co_i_1_7  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_8  co_1 co_i_1_8  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_9  co_1 co_i_1_9  VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_10 co_1 co_i_1_10 VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_11 co_1 co_i_1_11 VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_12 co_1 co_i_1_12 VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_13 co_1 co_i_1_13 VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_14 co_1 co_i_1_14 VGND int_con C=8f R=120
x_buf1_buf16_intcon_1_15 co_1 co_i_1_15 VGND int_con C=8f R=120

x16_0_0  co_i_0_0  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_0  sky130_fd_sc_hd__clkbuf_16
x16_0_1  co_i_0_1  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_1  sky130_fd_sc_hd__clkbuf_16
x16_0_2  co_i_0_2  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_2  sky130_fd_sc_hd__clkbuf_16
x16_0_3  co_i_0_3  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_3  sky130_fd_sc_hd__clkbuf_16
x16_0_4  co_i_0_4  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_4  sky130_fd_sc_hd__clkbuf_16
x16_0_5  co_i_0_5  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_5  sky130_fd_sc_hd__clkbuf_16
x16_0_6  co_i_0_6  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_6  sky130_fd_sc_hd__clkbuf_16
x16_0_7  co_i_0_7  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_7  sky130_fd_sc_hd__clkbuf_16
x16_0_8  co_i_0_8  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_8  sky130_fd_sc_hd__clkbuf_16
x16_0_9  co_i_0_9  VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_9  sky130_fd_sc_hd__clkbuf_16
x16_0_10 co_i_0_10 VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_10 sky130_fd_sc_hd__clkbuf_16
x16_0_11 co_i_0_11 VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_11 sky130_fd_sc_hd__clkbuf_16
x16_0_12 co_i_0_12 VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_12 sky130_fd_sc_hd__clkbuf_16
x16_0_13 co_i_0_13 VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_13 sky130_fd_sc_hd__clkbuf_16
x16_0_14 co_i_0_14 VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_14 sky130_fd_sc_hd__clkbuf_16
x16_0_15 co_i_0_15 VGND VNB vpwr_clk_buf1_0  vpwr_clk_buf1_0  ff_0_15 sky130_fd_sc_hd__clkbuf_16
x16_1_0  co_i_1_0  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_0  sky130_fd_sc_hd__clkbuf_16
x16_1_1  co_i_1_1  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_1  sky130_fd_sc_hd__clkbuf_16
x16_1_2  co_i_1_2  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_2  sky130_fd_sc_hd__clkbuf_16
x16_1_3  co_i_1_3  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_3  sky130_fd_sc_hd__clkbuf_16
x16_1_4  co_i_1_4  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_4  sky130_fd_sc_hd__clkbuf_16
x16_1_5  co_i_1_5  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_5  sky130_fd_sc_hd__clkbuf_16
x16_1_6  co_i_1_6  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_6  sky130_fd_sc_hd__clkbuf_16
x16_1_7  co_i_1_7  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_7  sky130_fd_sc_hd__clkbuf_16
x16_1_8  co_i_1_8  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_8  sky130_fd_sc_hd__clkbuf_16
x16_1_9  co_i_1_9  VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_9  sky130_fd_sc_hd__clkbuf_16
x16_1_10 co_i_1_10 VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_10 sky130_fd_sc_hd__clkbuf_16
x16_1_11 co_i_1_11 VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_11 sky130_fd_sc_hd__clkbuf_16
x16_1_12 co_i_1_12 VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_12 sky130_fd_sc_hd__clkbuf_16
x16_1_13 co_i_1_13 VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_13 sky130_fd_sc_hd__clkbuf_16
x16_1_14 co_i_1_14 VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_14 sky130_fd_sc_hd__clkbuf_16
x16_1_15 co_i_1_15 VGND VNB vpwr_clk_buf1_1  vpwr_clk_buf1_1  ff_1_15 sky130_fd_sc_hd__clkbuf_16

xf_0_0  ff_0_0  ff_clk_0_0  VGND ff_rc m=20
xf_0_1  ff_0_1  ff_clk_0_1  VGND ff_rc m=20
xf_0_2  ff_0_2  ff_clk_0_2  VGND ff_rc m=20
xf_0_3  ff_0_3  ff_clk_0_3  VGND ff_rc m=20
xf_0_4  ff_0_4  ff_clk_0_4  VGND ff_rc m=20
xf_0_5  ff_0_5  ff_clk_0_5  VGND ff_rc m=20
xf_0_6  ff_0_6  ff_clk_0_6  VGND ff_rc m=20
xf_0_7  ff_0_7  ff_clk_0_7  VGND ff_rc m=20
xf_0_8  ff_0_8  ff_clk_0_8  VGND ff_rc m=20
xf_0_9  ff_0_9  ff_clk_0_9  VGND ff_rc m=20
xf_0_10 ff_0_10 ff_clk_0_10 VGND ff_rc m=20
xf_0_11 ff_0_11 ff_clk_0_11 VGND ff_rc m=20
xf_0_12 ff_0_12 ff_clk_0_12 VGND ff_rc m=20
xf_0_13 ff_0_13 ff_clk_0_13 VGND ff_rc m=20
xf_0_14 ff_0_14 ff_clk_0_14 VGND ff_rc m=20
xf_0_15 ff_0_15 ff_clk_0_15 VGND ff_rc m=20
xf_1_0  ff_1_0  ff_clk_1_0  VGND ff_rc m=20
xf_1_1  ff_1_1  ff_clk_1_1  VGND ff_rc m=20
xf_1_2  ff_1_2  ff_clk_1_2  VGND ff_rc m=20
xf_1_3  ff_1_3  ff_clk_1_3  VGND ff_rc m=20
xf_1_4  ff_1_4  ff_clk_1_4  VGND ff_rc m=20
xf_1_5  ff_1_5  ff_clk_1_5  VGND ff_rc m=20
xf_1_6  ff_1_6  ff_clk_1_6  VGND ff_rc m=20
xf_1_7  ff_1_7  ff_clk_1_7  VGND ff_rc m=20
xf_1_8  ff_1_8  ff_clk_1_8  VGND ff_rc m=20
xf_1_9  ff_1_9  ff_clk_1_9  VGND ff_rc m=20
xf_1_10 ff_1_10 ff_clk_1_10 VGND ff_rc m=20
xf_1_11 ff_1_11 ff_clk_1_11 VGND ff_rc m=20
xf_1_12 ff_1_12 ff_clk_1_12 VGND ff_rc m=20
xf_1_13 ff_1_13 ff_clk_1_13 VGND ff_rc m=20
xf_1_14 ff_1_14 ff_clk_1_14 VGND ff_rc m=20
xf_1_15 ff_1_15 ff_clk_1_15 VGND ff_rc m=20

C_0_0 co_i_0_0  VGND 0.9F
C_0_1 co_i_0_1  VGND 0.9F
C_0_2 co_i_0_2  VGND 0.9F
C_0_3 co_i_0_3  VGND 0.9F
C_0_4 co_i_0_4  VGND 0.9F
C_0_5 co_i_0_5  VGND 0.9F
C_0_6 co_i_0_6  VGND 0.9F
C_0_7 co_i_0_7  VGND 0.9F
C_0_8 co_i_0_8  VGND 0.9F
C_0_9 co_i_0_9  VGND 0.9F
C_0_10 co_i_0_10 VGND 0.9F
C_0_11 co_i_0_11 VGND 0.9F
C_0_12 co_i_0_12 VGND 0.9F
C_0_13 co_i_0_13 VGND 0.9F
C_0_14 co_i_0_14 VGND 0.9F
C_0_15 co_i_0_15 VGND 0.9F
C_1_0 co_i_1_0  VGND 0.9F
C_1_1 co_i_1_1  VGND 0.9F
C_1_2 co_i_1_2  VGND 0.9F
C_1_3 co_i_1_3  VGND 0.9F
C_1_4 co_i_1_4  VGND 0.9F
C_1_5 co_i_1_5  VGND 0.9F
C_1_6 co_i_1_6  VGND 0.9F
C_1_7 co_i_1_7  VGND 0.9F
C_1_8 co_i_1_8  VGND 0.9F
C_1_9 co_i_1_9  VGND 0.9F
C_1_10 co_i_1_10 VGND 0.9F
C_1_11 co_i_1_11 VGND 0.9F
C_1_12 co_i_1_12 VGND 0.9F
C_1_13 co_i_1_13 VGND 0.9F
C_1_14 co_i_1_14 VGND 0.9F
C_1_15 co_i_1_15 VGND 0.9F


.lib     ../../../pdks/sky130A-1.0.227.01/libs.tech/ngspice/sky130.lib.spice tt
.include ../../../pdks/sky130A-1.0.227.01/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include ../../subckts.spice

.temp 25
.save all
.tran 0.1n 50n

.end

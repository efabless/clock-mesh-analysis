magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1515 -629 14693 6185
<< dnwell >>
rect 0 2004 12691 4841
rect 0 766 1205 2004
rect 4052 1954 12691 2004
rect 5461 766 12691 1954
<< nwell >>
rect -185 3937 13433 4925
rect -185 3629 10300 3937
rect -185 3615 84 3629
rect 897 3621 10300 3629
rect -255 3020 84 3615
rect 1948 3589 10300 3621
rect 1948 3476 3112 3589
rect -255 2164 32 3020
rect 12436 3341 13433 3937
rect 867 2164 1330 2240
rect -255 2024 1330 2164
rect 3110 2170 4530 2248
rect 3110 2070 5740 2170
rect 3110 2066 4530 2070
rect -255 1310 660 2024
rect -255 970 727 1310
rect 9089 1604 9287 2020
rect 10088 1713 10254 2335
rect 10146 1705 10254 1713
rect 12482 1705 13433 3341
rect 7971 970 8874 976
rect 12134 970 13433 1705
rect -255 631 13433 970
<< pwell >>
rect 9145 2873 9307 3525
rect 8437 1038 8727 1980
<< mvpsubdiff >>
rect 9171 3475 9281 3499
rect 9171 3441 9175 3475
rect 9209 3441 9243 3475
rect 9277 3441 9281 3475
rect 9171 3401 9281 3441
rect 9171 3367 9175 3401
rect 9209 3367 9243 3401
rect 9277 3367 9281 3401
rect 9171 3327 9281 3367
rect 9171 3293 9175 3327
rect 9209 3293 9243 3327
rect 9277 3293 9281 3327
rect 9171 3253 9281 3293
rect 9171 3219 9175 3253
rect 9209 3219 9243 3253
rect 9277 3219 9281 3253
rect 9171 3179 9281 3219
rect 9171 3145 9175 3179
rect 9209 3145 9243 3179
rect 9277 3145 9281 3179
rect 9171 3105 9281 3145
rect 9171 3071 9175 3105
rect 9209 3071 9243 3105
rect 9277 3071 9281 3105
rect 9171 3031 9281 3071
rect 9171 2997 9175 3031
rect 9209 2997 9243 3031
rect 9277 2997 9281 3031
rect 9171 2957 9281 2997
rect 9171 2923 9175 2957
rect 9209 2923 9243 2957
rect 9277 2923 9281 2957
rect 9171 2899 9281 2923
rect 8463 1930 8701 1954
rect 8497 1896 8531 1930
rect 8565 1896 8599 1930
rect 8633 1896 8667 1930
rect 8463 1856 8701 1896
rect 8497 1822 8531 1856
rect 8565 1822 8599 1856
rect 8633 1822 8667 1856
rect 8463 1782 8701 1822
rect 8497 1748 8531 1782
rect 8565 1748 8599 1782
rect 8633 1748 8667 1782
rect 8463 1708 8701 1748
rect 8497 1674 8531 1708
rect 8565 1674 8599 1708
rect 8633 1674 8667 1708
rect 8463 1634 8701 1674
rect 8497 1600 8531 1634
rect 8565 1600 8599 1634
rect 8633 1600 8667 1634
rect 8463 1560 8701 1600
rect 8497 1526 8531 1560
rect 8565 1526 8599 1560
rect 8633 1526 8667 1560
rect 8463 1487 8701 1526
rect 8497 1453 8531 1487
rect 8565 1453 8599 1487
rect 8633 1453 8667 1487
rect 8463 1414 8701 1453
rect 8497 1380 8531 1414
rect 8565 1380 8599 1414
rect 8633 1380 8667 1414
rect 8463 1341 8701 1380
rect 8497 1307 8531 1341
rect 8565 1307 8599 1341
rect 8633 1307 8667 1341
rect 8463 1268 8701 1307
rect 8497 1234 8531 1268
rect 8565 1234 8599 1268
rect 8633 1234 8667 1268
rect 8463 1195 8701 1234
rect 8497 1161 8531 1195
rect 8565 1161 8599 1195
rect 8633 1161 8667 1195
rect 8463 1122 8701 1161
rect 8497 1088 8531 1122
rect 8565 1088 8599 1122
rect 8633 1088 8667 1122
rect 8463 1064 8701 1088
<< mvnsubdiff >>
rect -17 4787 17 4858
rect 51 4824 161 4858
rect 195 4824 229 4858
rect 263 4824 297 4858
rect 331 4824 365 4858
rect 399 4824 433 4858
rect 467 4824 501 4858
rect 535 4824 569 4858
rect 603 4824 637 4858
rect 671 4824 705 4858
rect 739 4824 773 4858
rect 807 4824 841 4858
rect 875 4824 909 4858
rect 943 4824 977 4858
rect 1011 4824 1045 4858
rect 1079 4824 1113 4858
rect 1147 4824 1181 4858
rect 1215 4824 1249 4858
rect 1283 4824 1317 4858
rect 1351 4824 1385 4858
rect 1419 4824 1453 4858
rect 1487 4824 1521 4858
rect 1555 4824 1589 4858
rect 1623 4824 1657 4858
rect 1691 4824 1725 4858
rect 1759 4824 1793 4858
rect 1827 4824 1861 4858
rect 1895 4824 1929 4858
rect 1963 4824 1997 4858
rect 2031 4824 2065 4858
rect 2099 4824 2133 4858
rect 2167 4824 2201 4858
rect 2235 4824 2269 4858
rect 2303 4824 2337 4858
rect 2371 4824 2405 4858
rect 2439 4824 2473 4858
rect 2507 4824 2541 4858
rect 2575 4824 2609 4858
rect 2643 4824 2677 4858
rect 2711 4824 2745 4858
rect 2779 4824 2813 4858
rect 2847 4824 2881 4858
rect 2915 4824 2949 4858
rect 2983 4824 3017 4858
rect 3051 4824 3085 4858
rect 3119 4824 3153 4858
rect 3187 4824 3221 4858
rect 3255 4824 3289 4858
rect 3323 4824 3357 4858
rect 3391 4824 3425 4858
rect 3459 4824 3493 4858
rect 3527 4824 3561 4858
rect 3595 4824 3629 4858
rect 3663 4824 3697 4858
rect 3731 4824 3765 4858
rect 3799 4824 3833 4858
rect 3867 4824 3901 4858
rect 3935 4824 3969 4858
rect 4003 4824 4037 4858
rect 4071 4824 4105 4858
rect 4139 4824 4173 4858
rect 4207 4824 4241 4858
rect 4275 4824 4309 4858
rect 4343 4824 4377 4858
rect 4411 4824 4445 4858
rect 4479 4824 4513 4858
rect 4547 4824 4581 4858
rect 4615 4824 4649 4858
rect 4683 4824 4717 4858
rect 4751 4824 4785 4858
rect 4819 4824 4853 4858
rect 4887 4824 4921 4858
rect 4955 4824 4989 4858
rect 5023 4824 5057 4858
rect 5091 4824 5125 4858
rect 5159 4824 5193 4858
rect 5227 4824 5261 4858
rect 5295 4824 5329 4858
rect 5363 4824 5397 4858
rect 5431 4824 5465 4858
rect 5499 4824 5533 4858
rect 5567 4824 5601 4858
rect 5635 4824 5669 4858
rect 5703 4824 5737 4858
rect 5771 4824 5805 4858
rect 5839 4824 5873 4858
rect 5907 4824 5941 4858
rect 5975 4824 6009 4858
rect 6043 4824 6077 4858
rect 6111 4824 6145 4858
rect 6179 4824 6213 4858
rect 6247 4824 6281 4858
rect 6315 4824 6349 4858
rect 6383 4824 6417 4858
rect 6451 4824 6485 4858
rect 6519 4824 6553 4858
rect 6587 4824 6621 4858
rect 6655 4824 6689 4858
rect 6723 4824 6757 4858
rect 6791 4824 6825 4858
rect 6859 4824 6893 4858
rect 6927 4824 6961 4858
rect 6995 4824 7029 4858
rect 7063 4824 7097 4858
rect 7131 4824 7165 4858
rect 7199 4824 7233 4858
rect 7267 4824 7301 4858
rect 7335 4824 7369 4858
rect 7403 4824 7437 4858
rect 7471 4824 7505 4858
rect 7539 4824 7573 4858
rect 7607 4824 7641 4858
rect 7675 4824 7709 4858
rect 7743 4824 7777 4858
rect 7811 4824 7845 4858
rect 7879 4824 7913 4858
rect 7947 4824 7981 4858
rect 8015 4824 8049 4858
rect 8083 4824 8117 4858
rect 8151 4824 8185 4858
rect 8219 4824 8253 4858
rect 8287 4824 8321 4858
rect 8355 4824 8389 4858
rect 8423 4824 8457 4858
rect 8491 4824 8525 4858
rect 8559 4824 8593 4858
rect 8627 4824 8661 4858
rect 8695 4824 8729 4858
rect 8763 4824 8797 4858
rect 8831 4824 8865 4858
rect 8899 4824 8933 4858
rect 8967 4824 9001 4858
rect 9035 4824 9069 4858
rect 9103 4824 9137 4858
rect 9171 4824 9205 4858
rect 9239 4824 9273 4858
rect 9307 4824 9341 4858
rect 9375 4824 9409 4858
rect 9443 4824 9477 4858
rect 9511 4824 9545 4858
rect 9579 4824 9613 4858
rect 9647 4824 9681 4858
rect 9715 4824 9749 4858
rect 9783 4824 9817 4858
rect 9851 4824 9885 4858
rect 9919 4824 9953 4858
rect 9987 4824 10021 4858
rect 10055 4824 10089 4858
rect 10123 4824 10157 4858
rect 10191 4824 10225 4858
rect 10259 4824 10293 4858
rect 10327 4824 10361 4858
rect 10395 4824 10429 4858
rect 10463 4824 10497 4858
rect 10531 4824 10565 4858
rect 10599 4824 10633 4858
rect 10667 4824 10701 4858
rect 10735 4824 10769 4858
rect 10803 4824 10837 4858
rect 10871 4824 10905 4858
rect 10939 4824 10973 4858
rect 11007 4824 11041 4858
rect 11075 4824 11109 4858
rect 11143 4824 11177 4858
rect 11211 4824 11245 4858
rect 11279 4824 11313 4858
rect 11347 4824 11381 4858
rect 11415 4824 11449 4858
rect 11483 4824 11517 4858
rect 11551 4824 11585 4858
rect 11619 4824 11653 4858
rect 11687 4824 11721 4858
rect 11755 4824 11789 4858
rect 11823 4824 11857 4858
rect 11891 4824 11925 4858
rect 11959 4824 11993 4858
rect 12027 4824 12061 4858
rect 12095 4824 12129 4858
rect 12163 4824 12197 4858
rect 12231 4824 12265 4858
rect 12299 4824 12333 4858
rect 12367 4824 12401 4858
rect 12435 4824 12598 4858
rect -17 4719 17 4753
rect -17 4651 17 4685
rect -17 4583 17 4617
rect 12564 4758 12598 4824
rect 12564 4690 12598 4724
rect 12564 4622 12598 4656
rect -17 4515 17 4549
rect -17 4447 17 4481
rect -17 4379 17 4413
rect 321 4411 345 4581
rect 787 4411 811 4581
rect 12564 4554 12598 4588
rect 12564 4486 12598 4520
rect 12564 4418 12598 4452
rect -17 4311 17 4345
rect -17 4243 17 4277
rect -17 4175 17 4209
rect -17 4107 17 4141
rect -17 4039 17 4073
rect -17 3971 17 4005
rect -17 3903 17 3937
rect -17 3835 17 3869
rect 12564 4350 12598 4384
rect 12564 4282 12598 4316
rect 12564 4214 12598 4248
rect 12564 4146 12598 4180
rect 12564 4078 12598 4112
rect 12564 4010 12598 4044
rect 12564 3942 12598 3976
rect 12564 3874 12598 3908
rect -17 3767 17 3801
rect -17 3699 17 3733
rect -17 3631 17 3665
rect 10196 3655 10256 3825
rect 12564 3806 12598 3840
rect 12564 3738 12598 3772
rect 12564 3670 12598 3704
rect -17 3563 17 3597
rect -17 3495 17 3529
rect 12564 3602 12598 3636
rect 12564 3534 12598 3568
rect -17 3427 17 3461
rect -17 3359 17 3393
rect -17 3291 17 3325
rect -17 3223 17 3257
rect -17 3155 17 3189
rect -69 3087 17 3121
rect -69 3026 -35 3087
rect -69 2958 -35 2992
rect -69 2890 -35 2924
rect 12564 3466 12598 3500
rect 12564 3398 12598 3432
rect 12564 3330 12598 3364
rect 12564 3262 12598 3296
rect 12564 3194 12598 3228
rect 12564 3126 12598 3160
rect 12564 3058 12598 3092
rect 12564 2990 12598 3024
rect 12564 2922 12598 2956
rect -69 2822 -35 2856
rect -69 2754 -35 2788
rect -69 2686 -35 2720
rect -69 2618 -35 2652
rect -69 2550 -35 2584
rect -69 2482 -35 2516
rect -69 2414 -35 2448
rect -69 2346 -35 2380
rect -69 2278 -35 2312
rect 12564 2854 12598 2888
rect 12564 2786 12598 2820
rect 12564 2718 12598 2752
rect 12564 2650 12598 2684
rect 12564 2582 12598 2616
rect 12564 2514 12598 2548
rect 12564 2446 12598 2480
rect 12564 2378 12598 2412
rect 12564 2310 12598 2344
rect -69 2210 -35 2244
rect 10154 2245 10188 2269
rect -69 2142 -35 2176
rect 3176 2174 4464 2182
rect 3176 2140 3200 2174
rect 3234 2140 3271 2174
rect 3305 2140 3342 2174
rect 3376 2140 3413 2174
rect 3447 2140 3484 2174
rect 3518 2140 3555 2174
rect 3589 2140 3626 2174
rect 3660 2140 3697 2174
rect 3731 2140 3768 2174
rect 3802 2140 3839 2174
rect 3873 2140 3910 2174
rect 3944 2140 3981 2174
rect 4015 2140 4052 2174
rect 4086 2140 4123 2174
rect 4157 2140 4194 2174
rect 4228 2140 4265 2174
rect 4299 2140 4336 2174
rect 4370 2140 4406 2174
rect 4440 2140 4464 2174
rect 3176 2132 4464 2140
rect 10154 2177 10188 2211
rect -69 2074 -35 2108
rect -69 2006 -35 2040
rect -69 1938 -35 1972
rect 10154 2109 10188 2143
rect 10154 2041 10188 2075
rect 10154 1973 10188 2007
rect -69 1870 -35 1904
rect -69 1802 -35 1836
rect -69 1734 -35 1768
rect -69 1666 -35 1700
rect -69 1598 -35 1632
rect -69 1530 -35 1564
rect -69 1462 -35 1496
rect -69 1394 -35 1428
rect -69 1326 -35 1360
rect -69 1270 -35 1292
rect 9155 1930 9221 1954
rect 9155 1896 9171 1930
rect 9205 1896 9221 1930
rect 9155 1829 9221 1896
rect 9155 1795 9171 1829
rect 9205 1795 9221 1829
rect 9155 1728 9221 1795
rect 10154 1905 10188 1939
rect 10154 1837 10188 1871
rect 10154 1779 10188 1803
rect 12564 2242 12598 2276
rect 12564 2174 12598 2208
rect 12564 2106 12598 2140
rect 12564 2038 12598 2072
rect 12564 1970 12598 2004
rect 12564 1902 12598 1936
rect 12564 1834 12598 1868
rect 9155 1694 9171 1728
rect 9205 1694 9221 1728
rect 9155 1670 9221 1694
rect 12564 1766 12598 1800
rect 12564 1698 12598 1732
rect -69 1258 729 1270
rect -35 1224 729 1258
rect -69 1220 729 1224
rect -69 1190 83 1220
rect -35 1186 83 1190
rect 117 1186 151 1220
rect 185 1186 219 1220
rect 253 1186 287 1220
rect 321 1186 355 1220
rect 389 1186 423 1220
rect 457 1186 491 1220
rect 525 1186 559 1220
rect 593 1186 627 1220
rect 661 1186 729 1220
rect -35 1156 729 1186
rect -69 1151 729 1156
rect -69 1122 83 1151
rect -35 1117 83 1122
rect 117 1117 151 1151
rect 185 1117 219 1151
rect 253 1117 287 1151
rect 321 1117 355 1151
rect 389 1117 423 1151
rect 457 1117 491 1151
rect 525 1117 559 1151
rect 593 1117 627 1151
rect 661 1117 729 1151
rect -35 1088 729 1117
rect -69 1082 729 1088
rect -69 1054 83 1082
rect -35 1048 83 1054
rect 117 1048 151 1082
rect 185 1048 219 1082
rect 253 1048 287 1082
rect 321 1048 355 1082
rect 389 1048 423 1082
rect 457 1048 491 1082
rect 525 1048 559 1082
rect 593 1048 627 1082
rect 661 1048 729 1082
rect 12564 1630 12598 1664
rect 12564 1562 12598 1596
rect 12564 1494 12598 1528
rect 12564 1426 12598 1460
rect 12564 1358 12598 1392
rect 12564 1290 12598 1324
rect 12564 1222 12598 1256
rect 12564 1154 12598 1188
rect 12564 1086 12598 1120
rect -35 1020 729 1048
rect -69 1013 729 1020
rect -69 986 83 1013
rect -35 952 83 986
rect -69 918 83 952
rect -35 884 83 918
rect -69 850 83 884
rect -35 843 83 850
rect 661 843 729 1013
rect 12564 1018 12598 1052
rect 12564 950 12598 984
rect 12564 882 12598 916
rect 12564 846 12598 848
rect -35 816 729 843
rect -69 814 729 816
rect 12157 814 12598 846
rect -69 813 12564 814
rect -69 782 12190 813
rect -35 781 12190 782
rect -35 748 121 781
rect -69 747 121 748
rect 155 747 189 781
rect 223 747 257 781
rect 291 747 325 781
rect 359 747 393 781
rect 427 747 461 781
rect 495 747 529 781
rect 563 747 597 781
rect 631 747 665 781
rect 699 747 733 781
rect 767 747 801 781
rect 835 747 869 781
rect 903 747 937 781
rect 971 747 1005 781
rect 1039 747 1073 781
rect 1107 747 1141 781
rect 1175 747 1209 781
rect 1243 747 1277 781
rect 1311 747 1345 781
rect 1379 747 1413 781
rect 1447 747 1481 781
rect 1515 747 1549 781
rect 1583 747 1617 781
rect 1651 747 1685 781
rect 1719 747 1753 781
rect 1787 747 1821 781
rect 1855 747 1889 781
rect 1923 747 1957 781
rect 1991 747 2025 781
rect 2059 747 2093 781
rect 2127 747 2161 781
rect 2195 747 2229 781
rect 2263 747 2297 781
rect 2331 747 2365 781
rect 2399 747 2433 781
rect 2467 747 2501 781
rect 2535 747 2569 781
rect 2603 747 2637 781
rect 2671 747 2705 781
rect 2739 747 2773 781
rect 2807 747 2841 781
rect 2875 747 2909 781
rect 2943 747 2977 781
rect 3011 747 3045 781
rect 3079 747 3113 781
rect 3147 747 3181 781
rect 3215 747 3249 781
rect 3283 747 3317 781
rect 3351 747 3385 781
rect 3419 747 3453 781
rect 3487 747 3521 781
rect 3555 747 3589 781
rect 3623 747 3657 781
rect 3691 747 3725 781
rect 3759 747 3793 781
rect 3827 747 3861 781
rect 3895 747 3929 781
rect 3963 747 3997 781
rect 4031 747 4065 781
rect 4099 747 4133 781
rect 4167 747 4201 781
rect 4235 747 4269 781
rect 4303 747 4337 781
rect 4371 747 4405 781
rect 4439 747 4473 781
rect 4507 747 4541 781
rect 4575 747 4609 781
rect 4643 747 4677 781
rect 4711 747 4745 781
rect 4779 747 4813 781
rect 4847 747 4881 781
rect 4915 747 4949 781
rect 4983 747 5017 781
rect 5051 747 5085 781
rect 5119 747 5153 781
rect 5187 747 5221 781
rect 5255 747 5289 781
rect 5323 747 5357 781
rect 5391 747 5425 781
rect 5459 747 5493 781
rect 5527 747 5561 781
rect 5595 747 5629 781
rect 5663 747 5697 781
rect 5731 747 5765 781
rect 5799 747 5833 781
rect 5867 747 5901 781
rect 5935 747 5969 781
rect 6003 747 6037 781
rect 6071 747 6105 781
rect 6139 747 6173 781
rect 6207 747 6241 781
rect 6275 747 6309 781
rect 6343 747 6377 781
rect 6411 747 6445 781
rect 6479 747 6513 781
rect 6547 747 6581 781
rect 6615 747 6649 781
rect 6683 747 6717 781
rect 6751 747 6785 781
rect 6819 747 6853 781
rect 6887 747 6921 781
rect 6955 747 6989 781
rect 7023 747 7057 781
rect 7091 747 7125 781
rect 7159 747 7193 781
rect 7227 747 7261 781
rect 7295 747 7329 781
rect 7363 747 7397 781
rect 7431 747 7465 781
rect 7499 747 7533 781
rect 7567 747 7601 781
rect 7635 747 7669 781
rect 7703 747 7737 781
rect 7771 747 7805 781
rect 7839 747 7873 781
rect 7907 747 7941 781
rect 7975 747 8009 781
rect 8043 747 8077 781
rect 8111 747 8145 781
rect 8179 747 8213 781
rect 8247 747 8281 781
rect 8315 747 8349 781
rect 8383 747 8417 781
rect 8451 747 8485 781
rect 8519 747 8553 781
rect 8587 747 8621 781
rect 8655 747 8689 781
rect 8723 747 8757 781
rect 8791 747 8825 781
rect 8859 747 8893 781
rect 8927 747 8961 781
rect 8995 747 9029 781
rect 9063 747 9097 781
rect 9131 747 9165 781
rect 9199 747 9233 781
rect 9267 747 9301 781
rect 9335 747 9369 781
rect 9403 747 9437 781
rect 9471 747 9505 781
rect 9539 747 9573 781
rect 9607 747 9641 781
rect 9675 747 9709 781
rect 9743 747 9777 781
rect 9811 747 9845 781
rect 9879 747 9913 781
rect 9947 747 9981 781
rect 10015 747 10049 781
rect 10083 747 10117 781
rect 10151 747 10185 781
rect 10219 747 10253 781
rect 10287 747 10321 781
rect 10355 747 10389 781
rect 10423 747 10457 781
rect 10491 747 10525 781
rect 10559 747 10593 781
rect 10627 747 10661 781
rect 10695 747 10729 781
rect 10763 747 10797 781
rect 10831 747 10865 781
rect 10899 747 10933 781
rect 10967 747 11001 781
rect 11035 747 11069 781
rect 11103 747 11137 781
rect 11171 747 11205 781
rect 11239 747 11273 781
rect 11307 747 11341 781
rect 11375 747 11409 781
rect 11443 747 11477 781
rect 11511 747 11545 781
rect 11579 747 11613 781
rect 11647 747 11681 781
rect 11715 747 11749 781
rect 11783 747 11817 781
rect 11851 747 11885 781
rect 11919 747 11953 781
rect 11987 747 12021 781
rect 12055 747 12089 781
rect 12123 779 12190 781
rect 12224 779 12258 813
rect 12292 779 12326 813
rect 12360 779 12394 813
rect 12428 779 12462 813
rect 12496 780 12564 813
rect 12496 779 12598 780
rect 12123 747 12598 779
rect -69 746 12598 747
rect -69 714 12257 746
<< mvpsubdiffcont >>
rect 9175 3441 9209 3475
rect 9243 3441 9277 3475
rect 9175 3367 9209 3401
rect 9243 3367 9277 3401
rect 9175 3293 9209 3327
rect 9243 3293 9277 3327
rect 9175 3219 9209 3253
rect 9243 3219 9277 3253
rect 9175 3145 9209 3179
rect 9243 3145 9277 3179
rect 9175 3071 9209 3105
rect 9243 3071 9277 3105
rect 9175 2997 9209 3031
rect 9243 2997 9277 3031
rect 9175 2923 9209 2957
rect 9243 2923 9277 2957
rect 8463 1896 8497 1930
rect 8531 1896 8565 1930
rect 8599 1896 8633 1930
rect 8667 1896 8701 1930
rect 8463 1822 8497 1856
rect 8531 1822 8565 1856
rect 8599 1822 8633 1856
rect 8667 1822 8701 1856
rect 8463 1748 8497 1782
rect 8531 1748 8565 1782
rect 8599 1748 8633 1782
rect 8667 1748 8701 1782
rect 8463 1674 8497 1708
rect 8531 1674 8565 1708
rect 8599 1674 8633 1708
rect 8667 1674 8701 1708
rect 8463 1600 8497 1634
rect 8531 1600 8565 1634
rect 8599 1600 8633 1634
rect 8667 1600 8701 1634
rect 8463 1526 8497 1560
rect 8531 1526 8565 1560
rect 8599 1526 8633 1560
rect 8667 1526 8701 1560
rect 8463 1453 8497 1487
rect 8531 1453 8565 1487
rect 8599 1453 8633 1487
rect 8667 1453 8701 1487
rect 8463 1380 8497 1414
rect 8531 1380 8565 1414
rect 8599 1380 8633 1414
rect 8667 1380 8701 1414
rect 8463 1307 8497 1341
rect 8531 1307 8565 1341
rect 8599 1307 8633 1341
rect 8667 1307 8701 1341
rect 8463 1234 8497 1268
rect 8531 1234 8565 1268
rect 8599 1234 8633 1268
rect 8667 1234 8701 1268
rect 8463 1161 8497 1195
rect 8531 1161 8565 1195
rect 8599 1161 8633 1195
rect 8667 1161 8701 1195
rect 8463 1088 8497 1122
rect 8531 1088 8565 1122
rect 8599 1088 8633 1122
rect 8667 1088 8701 1122
<< mvnsubdiffcont >>
rect 17 4824 51 4858
rect 161 4824 195 4858
rect 229 4824 263 4858
rect 297 4824 331 4858
rect 365 4824 399 4858
rect 433 4824 467 4858
rect 501 4824 535 4858
rect 569 4824 603 4858
rect 637 4824 671 4858
rect 705 4824 739 4858
rect 773 4824 807 4858
rect 841 4824 875 4858
rect 909 4824 943 4858
rect 977 4824 1011 4858
rect 1045 4824 1079 4858
rect 1113 4824 1147 4858
rect 1181 4824 1215 4858
rect 1249 4824 1283 4858
rect 1317 4824 1351 4858
rect 1385 4824 1419 4858
rect 1453 4824 1487 4858
rect 1521 4824 1555 4858
rect 1589 4824 1623 4858
rect 1657 4824 1691 4858
rect 1725 4824 1759 4858
rect 1793 4824 1827 4858
rect 1861 4824 1895 4858
rect 1929 4824 1963 4858
rect 1997 4824 2031 4858
rect 2065 4824 2099 4858
rect 2133 4824 2167 4858
rect 2201 4824 2235 4858
rect 2269 4824 2303 4858
rect 2337 4824 2371 4858
rect 2405 4824 2439 4858
rect 2473 4824 2507 4858
rect 2541 4824 2575 4858
rect 2609 4824 2643 4858
rect 2677 4824 2711 4858
rect 2745 4824 2779 4858
rect 2813 4824 2847 4858
rect 2881 4824 2915 4858
rect 2949 4824 2983 4858
rect 3017 4824 3051 4858
rect 3085 4824 3119 4858
rect 3153 4824 3187 4858
rect 3221 4824 3255 4858
rect 3289 4824 3323 4858
rect 3357 4824 3391 4858
rect 3425 4824 3459 4858
rect 3493 4824 3527 4858
rect 3561 4824 3595 4858
rect 3629 4824 3663 4858
rect 3697 4824 3731 4858
rect 3765 4824 3799 4858
rect 3833 4824 3867 4858
rect 3901 4824 3935 4858
rect 3969 4824 4003 4858
rect 4037 4824 4071 4858
rect 4105 4824 4139 4858
rect 4173 4824 4207 4858
rect 4241 4824 4275 4858
rect 4309 4824 4343 4858
rect 4377 4824 4411 4858
rect 4445 4824 4479 4858
rect 4513 4824 4547 4858
rect 4581 4824 4615 4858
rect 4649 4824 4683 4858
rect 4717 4824 4751 4858
rect 4785 4824 4819 4858
rect 4853 4824 4887 4858
rect 4921 4824 4955 4858
rect 4989 4824 5023 4858
rect 5057 4824 5091 4858
rect 5125 4824 5159 4858
rect 5193 4824 5227 4858
rect 5261 4824 5295 4858
rect 5329 4824 5363 4858
rect 5397 4824 5431 4858
rect 5465 4824 5499 4858
rect 5533 4824 5567 4858
rect 5601 4824 5635 4858
rect 5669 4824 5703 4858
rect 5737 4824 5771 4858
rect 5805 4824 5839 4858
rect 5873 4824 5907 4858
rect 5941 4824 5975 4858
rect 6009 4824 6043 4858
rect 6077 4824 6111 4858
rect 6145 4824 6179 4858
rect 6213 4824 6247 4858
rect 6281 4824 6315 4858
rect 6349 4824 6383 4858
rect 6417 4824 6451 4858
rect 6485 4824 6519 4858
rect 6553 4824 6587 4858
rect 6621 4824 6655 4858
rect 6689 4824 6723 4858
rect 6757 4824 6791 4858
rect 6825 4824 6859 4858
rect 6893 4824 6927 4858
rect 6961 4824 6995 4858
rect 7029 4824 7063 4858
rect 7097 4824 7131 4858
rect 7165 4824 7199 4858
rect 7233 4824 7267 4858
rect 7301 4824 7335 4858
rect 7369 4824 7403 4858
rect 7437 4824 7471 4858
rect 7505 4824 7539 4858
rect 7573 4824 7607 4858
rect 7641 4824 7675 4858
rect 7709 4824 7743 4858
rect 7777 4824 7811 4858
rect 7845 4824 7879 4858
rect 7913 4824 7947 4858
rect 7981 4824 8015 4858
rect 8049 4824 8083 4858
rect 8117 4824 8151 4858
rect 8185 4824 8219 4858
rect 8253 4824 8287 4858
rect 8321 4824 8355 4858
rect 8389 4824 8423 4858
rect 8457 4824 8491 4858
rect 8525 4824 8559 4858
rect 8593 4824 8627 4858
rect 8661 4824 8695 4858
rect 8729 4824 8763 4858
rect 8797 4824 8831 4858
rect 8865 4824 8899 4858
rect 8933 4824 8967 4858
rect 9001 4824 9035 4858
rect 9069 4824 9103 4858
rect 9137 4824 9171 4858
rect 9205 4824 9239 4858
rect 9273 4824 9307 4858
rect 9341 4824 9375 4858
rect 9409 4824 9443 4858
rect 9477 4824 9511 4858
rect 9545 4824 9579 4858
rect 9613 4824 9647 4858
rect 9681 4824 9715 4858
rect 9749 4824 9783 4858
rect 9817 4824 9851 4858
rect 9885 4824 9919 4858
rect 9953 4824 9987 4858
rect 10021 4824 10055 4858
rect 10089 4824 10123 4858
rect 10157 4824 10191 4858
rect 10225 4824 10259 4858
rect 10293 4824 10327 4858
rect 10361 4824 10395 4858
rect 10429 4824 10463 4858
rect 10497 4824 10531 4858
rect 10565 4824 10599 4858
rect 10633 4824 10667 4858
rect 10701 4824 10735 4858
rect 10769 4824 10803 4858
rect 10837 4824 10871 4858
rect 10905 4824 10939 4858
rect 10973 4824 11007 4858
rect 11041 4824 11075 4858
rect 11109 4824 11143 4858
rect 11177 4824 11211 4858
rect 11245 4824 11279 4858
rect 11313 4824 11347 4858
rect 11381 4824 11415 4858
rect 11449 4824 11483 4858
rect 11517 4824 11551 4858
rect 11585 4824 11619 4858
rect 11653 4824 11687 4858
rect 11721 4824 11755 4858
rect 11789 4824 11823 4858
rect 11857 4824 11891 4858
rect 11925 4824 11959 4858
rect 11993 4824 12027 4858
rect 12061 4824 12095 4858
rect 12129 4824 12163 4858
rect 12197 4824 12231 4858
rect 12265 4824 12299 4858
rect 12333 4824 12367 4858
rect 12401 4824 12435 4858
rect -17 4753 17 4787
rect -17 4685 17 4719
rect -17 4617 17 4651
rect -17 4549 17 4583
rect 12564 4724 12598 4758
rect 12564 4656 12598 4690
rect 12564 4588 12598 4622
rect -17 4481 17 4515
rect -17 4413 17 4447
rect 345 4411 787 4581
rect 12564 4520 12598 4554
rect 12564 4452 12598 4486
rect -17 4345 17 4379
rect -17 4277 17 4311
rect -17 4209 17 4243
rect -17 4141 17 4175
rect -17 4073 17 4107
rect -17 4005 17 4039
rect -17 3937 17 3971
rect -17 3869 17 3903
rect -17 3801 17 3835
rect 12564 4384 12598 4418
rect 12564 4316 12598 4350
rect 12564 4248 12598 4282
rect 12564 4180 12598 4214
rect 12564 4112 12598 4146
rect 12564 4044 12598 4078
rect 12564 3976 12598 4010
rect 12564 3908 12598 3942
rect 12564 3840 12598 3874
rect -17 3733 17 3767
rect -17 3665 17 3699
rect 12564 3772 12598 3806
rect 12564 3704 12598 3738
rect -17 3597 17 3631
rect -17 3529 17 3563
rect 12564 3636 12598 3670
rect 12564 3568 12598 3602
rect 12564 3500 12598 3534
rect -17 3461 17 3495
rect -17 3393 17 3427
rect -17 3325 17 3359
rect -17 3257 17 3291
rect -17 3189 17 3223
rect -17 3121 17 3155
rect -69 2992 -35 3026
rect -69 2924 -35 2958
rect 12564 3432 12598 3466
rect 12564 3364 12598 3398
rect 12564 3296 12598 3330
rect 12564 3228 12598 3262
rect 12564 3160 12598 3194
rect 12564 3092 12598 3126
rect 12564 3024 12598 3058
rect 12564 2956 12598 2990
rect -69 2856 -35 2890
rect -69 2788 -35 2822
rect -69 2720 -35 2754
rect -69 2652 -35 2686
rect -69 2584 -35 2618
rect -69 2516 -35 2550
rect -69 2448 -35 2482
rect -69 2380 -35 2414
rect -69 2312 -35 2346
rect -69 2244 -35 2278
rect 12564 2888 12598 2922
rect 12564 2820 12598 2854
rect 12564 2752 12598 2786
rect 12564 2684 12598 2718
rect 12564 2616 12598 2650
rect 12564 2548 12598 2582
rect 12564 2480 12598 2514
rect 12564 2412 12598 2446
rect 12564 2344 12598 2378
rect 12564 2276 12598 2310
rect -69 2176 -35 2210
rect 10154 2211 10188 2245
rect -69 2108 -35 2142
rect 3200 2140 3234 2174
rect 3271 2140 3305 2174
rect 3342 2140 3376 2174
rect 3413 2140 3447 2174
rect 3484 2140 3518 2174
rect 3555 2140 3589 2174
rect 3626 2140 3660 2174
rect 3697 2140 3731 2174
rect 3768 2140 3802 2174
rect 3839 2140 3873 2174
rect 3910 2140 3944 2174
rect 3981 2140 4015 2174
rect 4052 2140 4086 2174
rect 4123 2140 4157 2174
rect 4194 2140 4228 2174
rect 4265 2140 4299 2174
rect 4336 2140 4370 2174
rect 4406 2140 4440 2174
rect 10154 2143 10188 2177
rect -69 2040 -35 2074
rect -69 1972 -35 2006
rect 10154 2075 10188 2109
rect 10154 2007 10188 2041
rect -69 1904 -35 1938
rect -69 1836 -35 1870
rect -69 1768 -35 1802
rect -69 1700 -35 1734
rect -69 1632 -35 1666
rect -69 1564 -35 1598
rect -69 1496 -35 1530
rect -69 1428 -35 1462
rect -69 1360 -35 1394
rect -69 1292 -35 1326
rect 9171 1896 9205 1930
rect 9171 1795 9205 1829
rect 10154 1939 10188 1973
rect 10154 1871 10188 1905
rect 10154 1803 10188 1837
rect 12564 2208 12598 2242
rect 12564 2140 12598 2174
rect 12564 2072 12598 2106
rect 12564 2004 12598 2038
rect 12564 1936 12598 1970
rect 12564 1868 12598 1902
rect 12564 1800 12598 1834
rect 9171 1694 9205 1728
rect 12564 1732 12598 1766
rect -69 1224 -35 1258
rect -69 1156 -35 1190
rect 83 1186 117 1220
rect 151 1186 185 1220
rect 219 1186 253 1220
rect 287 1186 321 1220
rect 355 1186 389 1220
rect 423 1186 457 1220
rect 491 1186 525 1220
rect 559 1186 593 1220
rect 627 1186 661 1220
rect -69 1088 -35 1122
rect 83 1117 117 1151
rect 151 1117 185 1151
rect 219 1117 253 1151
rect 287 1117 321 1151
rect 355 1117 389 1151
rect 423 1117 457 1151
rect 491 1117 525 1151
rect 559 1117 593 1151
rect 627 1117 661 1151
rect -69 1020 -35 1054
rect 83 1048 117 1082
rect 151 1048 185 1082
rect 219 1048 253 1082
rect 287 1048 321 1082
rect 355 1048 389 1082
rect 423 1048 457 1082
rect 491 1048 525 1082
rect 559 1048 593 1082
rect 627 1048 661 1082
rect 12564 1664 12598 1698
rect 12564 1596 12598 1630
rect 12564 1528 12598 1562
rect 12564 1460 12598 1494
rect 12564 1392 12598 1426
rect 12564 1324 12598 1358
rect 12564 1256 12598 1290
rect 12564 1188 12598 1222
rect 12564 1120 12598 1154
rect -69 952 -35 986
rect -69 884 -35 918
rect -69 816 -35 850
rect 83 843 661 1013
rect 12564 1052 12598 1086
rect 12564 984 12598 1018
rect 12564 916 12598 950
rect 12564 848 12598 882
rect -69 748 -35 782
rect 121 747 155 781
rect 189 747 223 781
rect 257 747 291 781
rect 325 747 359 781
rect 393 747 427 781
rect 461 747 495 781
rect 529 747 563 781
rect 597 747 631 781
rect 665 747 699 781
rect 733 747 767 781
rect 801 747 835 781
rect 869 747 903 781
rect 937 747 971 781
rect 1005 747 1039 781
rect 1073 747 1107 781
rect 1141 747 1175 781
rect 1209 747 1243 781
rect 1277 747 1311 781
rect 1345 747 1379 781
rect 1413 747 1447 781
rect 1481 747 1515 781
rect 1549 747 1583 781
rect 1617 747 1651 781
rect 1685 747 1719 781
rect 1753 747 1787 781
rect 1821 747 1855 781
rect 1889 747 1923 781
rect 1957 747 1991 781
rect 2025 747 2059 781
rect 2093 747 2127 781
rect 2161 747 2195 781
rect 2229 747 2263 781
rect 2297 747 2331 781
rect 2365 747 2399 781
rect 2433 747 2467 781
rect 2501 747 2535 781
rect 2569 747 2603 781
rect 2637 747 2671 781
rect 2705 747 2739 781
rect 2773 747 2807 781
rect 2841 747 2875 781
rect 2909 747 2943 781
rect 2977 747 3011 781
rect 3045 747 3079 781
rect 3113 747 3147 781
rect 3181 747 3215 781
rect 3249 747 3283 781
rect 3317 747 3351 781
rect 3385 747 3419 781
rect 3453 747 3487 781
rect 3521 747 3555 781
rect 3589 747 3623 781
rect 3657 747 3691 781
rect 3725 747 3759 781
rect 3793 747 3827 781
rect 3861 747 3895 781
rect 3929 747 3963 781
rect 3997 747 4031 781
rect 4065 747 4099 781
rect 4133 747 4167 781
rect 4201 747 4235 781
rect 4269 747 4303 781
rect 4337 747 4371 781
rect 4405 747 4439 781
rect 4473 747 4507 781
rect 4541 747 4575 781
rect 4609 747 4643 781
rect 4677 747 4711 781
rect 4745 747 4779 781
rect 4813 747 4847 781
rect 4881 747 4915 781
rect 4949 747 4983 781
rect 5017 747 5051 781
rect 5085 747 5119 781
rect 5153 747 5187 781
rect 5221 747 5255 781
rect 5289 747 5323 781
rect 5357 747 5391 781
rect 5425 747 5459 781
rect 5493 747 5527 781
rect 5561 747 5595 781
rect 5629 747 5663 781
rect 5697 747 5731 781
rect 5765 747 5799 781
rect 5833 747 5867 781
rect 5901 747 5935 781
rect 5969 747 6003 781
rect 6037 747 6071 781
rect 6105 747 6139 781
rect 6173 747 6207 781
rect 6241 747 6275 781
rect 6309 747 6343 781
rect 6377 747 6411 781
rect 6445 747 6479 781
rect 6513 747 6547 781
rect 6581 747 6615 781
rect 6649 747 6683 781
rect 6717 747 6751 781
rect 6785 747 6819 781
rect 6853 747 6887 781
rect 6921 747 6955 781
rect 6989 747 7023 781
rect 7057 747 7091 781
rect 7125 747 7159 781
rect 7193 747 7227 781
rect 7261 747 7295 781
rect 7329 747 7363 781
rect 7397 747 7431 781
rect 7465 747 7499 781
rect 7533 747 7567 781
rect 7601 747 7635 781
rect 7669 747 7703 781
rect 7737 747 7771 781
rect 7805 747 7839 781
rect 7873 747 7907 781
rect 7941 747 7975 781
rect 8009 747 8043 781
rect 8077 747 8111 781
rect 8145 747 8179 781
rect 8213 747 8247 781
rect 8281 747 8315 781
rect 8349 747 8383 781
rect 8417 747 8451 781
rect 8485 747 8519 781
rect 8553 747 8587 781
rect 8621 747 8655 781
rect 8689 747 8723 781
rect 8757 747 8791 781
rect 8825 747 8859 781
rect 8893 747 8927 781
rect 8961 747 8995 781
rect 9029 747 9063 781
rect 9097 747 9131 781
rect 9165 747 9199 781
rect 9233 747 9267 781
rect 9301 747 9335 781
rect 9369 747 9403 781
rect 9437 747 9471 781
rect 9505 747 9539 781
rect 9573 747 9607 781
rect 9641 747 9675 781
rect 9709 747 9743 781
rect 9777 747 9811 781
rect 9845 747 9879 781
rect 9913 747 9947 781
rect 9981 747 10015 781
rect 10049 747 10083 781
rect 10117 747 10151 781
rect 10185 747 10219 781
rect 10253 747 10287 781
rect 10321 747 10355 781
rect 10389 747 10423 781
rect 10457 747 10491 781
rect 10525 747 10559 781
rect 10593 747 10627 781
rect 10661 747 10695 781
rect 10729 747 10763 781
rect 10797 747 10831 781
rect 10865 747 10899 781
rect 10933 747 10967 781
rect 11001 747 11035 781
rect 11069 747 11103 781
rect 11137 747 11171 781
rect 11205 747 11239 781
rect 11273 747 11307 781
rect 11341 747 11375 781
rect 11409 747 11443 781
rect 11477 747 11511 781
rect 11545 747 11579 781
rect 11613 747 11647 781
rect 11681 747 11715 781
rect 11749 747 11783 781
rect 11817 747 11851 781
rect 11885 747 11919 781
rect 11953 747 11987 781
rect 12021 747 12055 781
rect 12089 747 12123 781
rect 12190 779 12224 813
rect 12258 779 12292 813
rect 12326 779 12360 813
rect 12394 779 12428 813
rect 12462 779 12496 813
rect 12564 780 12598 814
<< locali >>
rect 51 4824 55 4858
rect 89 4824 127 4858
rect 195 4824 199 4858
rect 263 4824 271 4858
rect 331 4824 343 4858
rect 399 4824 415 4858
rect 467 4824 501 4858
rect 542 4824 569 4858
rect 614 4824 637 4858
rect 686 4824 705 4858
rect 758 4824 773 4858
rect 830 4824 841 4858
rect 902 4824 909 4858
rect 974 4824 977 4858
rect 1011 4824 1012 4858
rect 1079 4824 1084 4858
rect 1147 4824 1156 4858
rect 1215 4824 1228 4858
rect 1283 4824 1300 4858
rect 1351 4824 1372 4858
rect 1419 4824 1444 4858
rect 1487 4824 1516 4858
rect 1555 4824 1588 4858
rect 1623 4824 1657 4858
rect 1694 4824 1725 4858
rect 1766 4824 1793 4858
rect 1838 4824 1861 4858
rect 1910 4824 1929 4858
rect 1982 4824 1997 4858
rect 2054 4824 2065 4858
rect 2126 4824 2133 4858
rect 2198 4824 2201 4858
rect 2235 4824 2236 4858
rect 2303 4824 2308 4858
rect 2371 4824 2380 4858
rect 2439 4824 2452 4858
rect 2507 4824 2524 4858
rect 2575 4824 2596 4858
rect 2643 4824 2668 4858
rect 2711 4824 2740 4858
rect 2779 4824 2812 4858
rect 2847 4824 2881 4858
rect 2918 4824 2949 4858
rect 2990 4824 3017 4858
rect 3062 4824 3085 4858
rect 3134 4824 3153 4858
rect 3206 4824 3221 4858
rect 3278 4824 3289 4858
rect 3350 4824 3357 4858
rect 3422 4824 3425 4858
rect 3459 4824 3460 4858
rect 3527 4824 3532 4858
rect 3595 4824 3604 4858
rect 3663 4824 3676 4858
rect 3731 4824 3748 4858
rect 3799 4824 3820 4858
rect 3867 4824 3892 4858
rect 3935 4824 3964 4858
rect 4003 4824 4036 4858
rect 4071 4824 4105 4858
rect 4142 4824 4173 4858
rect 4214 4824 4241 4858
rect 4286 4824 4309 4858
rect 4358 4824 4377 4858
rect 4430 4824 4445 4858
rect 4502 4824 4513 4858
rect 4574 4824 4581 4858
rect 4646 4824 4649 4858
rect 4683 4824 4684 4858
rect 4751 4824 4756 4858
rect 4819 4824 4828 4858
rect 4887 4824 4900 4858
rect 4955 4824 4972 4858
rect 5023 4824 5044 4858
rect 5091 4824 5116 4858
rect 5159 4824 5188 4858
rect 5227 4824 5260 4858
rect 5295 4824 5329 4858
rect 5366 4824 5397 4858
rect 5438 4824 5465 4858
rect 5510 4824 5533 4858
rect 5582 4824 5601 4858
rect 5654 4824 5669 4858
rect 5726 4824 5737 4858
rect 5798 4824 5805 4858
rect 5870 4824 5873 4858
rect 5907 4824 5908 4858
rect 5975 4824 5980 4858
rect 6043 4824 6052 4858
rect 6111 4824 6124 4858
rect 6179 4824 6196 4858
rect 6247 4824 6268 4858
rect 6315 4824 6340 4858
rect 6383 4824 6412 4858
rect 6451 4824 6484 4858
rect 6519 4824 6553 4858
rect 6590 4824 6621 4858
rect 6662 4824 6689 4858
rect 6734 4824 6757 4858
rect 6806 4824 6825 4858
rect 6878 4824 6893 4858
rect 6950 4824 6961 4858
rect 7022 4824 7029 4858
rect 7094 4824 7097 4858
rect 7131 4824 7132 4858
rect 7199 4824 7204 4858
rect 7267 4824 7276 4858
rect 7335 4824 7348 4858
rect 7403 4824 7420 4858
rect 7471 4824 7492 4858
rect 7539 4824 7564 4858
rect 7607 4824 7636 4858
rect 7675 4824 7708 4858
rect 7743 4824 7777 4858
rect 7814 4824 7845 4858
rect 7886 4824 7913 4858
rect 7958 4824 7981 4858
rect 8030 4824 8049 4858
rect 8102 4824 8117 4858
rect 8174 4824 8185 4858
rect 8246 4824 8253 4858
rect 8318 4824 8321 4858
rect 8355 4824 8356 4858
rect 8423 4824 8428 4858
rect 8491 4824 8500 4858
rect 8559 4824 8572 4858
rect 8627 4824 8644 4858
rect 8695 4824 8716 4858
rect 8763 4824 8788 4858
rect 8831 4824 8860 4858
rect 8899 4824 8932 4858
rect 8967 4824 9001 4858
rect 9038 4824 9069 4858
rect 9110 4824 9137 4858
rect 9182 4824 9205 4858
rect 9254 4824 9273 4858
rect 9326 4824 9341 4858
rect 9398 4824 9409 4858
rect 9470 4824 9477 4858
rect 9542 4824 9545 4858
rect 9579 4824 9580 4858
rect 9647 4824 9652 4858
rect 9715 4824 9724 4858
rect 9783 4824 9796 4858
rect 9851 4824 9868 4858
rect 9919 4824 9940 4858
rect 9987 4824 10012 4858
rect 10055 4824 10084 4858
rect 10123 4824 10156 4858
rect 10191 4824 10225 4858
rect 10262 4824 10293 4858
rect 10334 4824 10361 4858
rect 10406 4824 10429 4858
rect 10478 4824 10497 4858
rect 10550 4824 10565 4858
rect 10622 4824 10633 4858
rect 10694 4824 10701 4858
rect 10766 4824 10769 4858
rect 10803 4824 10804 4858
rect 10871 4824 10876 4858
rect 10939 4824 10948 4858
rect 11007 4824 11020 4858
rect 11075 4824 11092 4858
rect 11143 4824 11164 4858
rect 11211 4824 11236 4858
rect 11279 4824 11308 4858
rect 11347 4824 11380 4858
rect 11415 4824 11449 4858
rect 11486 4824 11517 4858
rect 11558 4824 11585 4858
rect 11630 4824 11653 4858
rect 11702 4824 11721 4858
rect 11774 4824 11789 4858
rect 11847 4824 11857 4858
rect 11920 4824 11925 4858
rect 12027 4824 12032 4858
rect 12095 4824 12105 4858
rect 12163 4824 12178 4858
rect 12231 4824 12251 4858
rect 12299 4824 12324 4858
rect 12367 4824 12397 4858
rect 12435 4824 12470 4858
rect 12504 4824 12543 4858
rect 12577 4824 12616 4858
rect 12650 4824 12689 4858
rect 12723 4824 12762 4858
rect 12796 4824 12835 4858
rect 12869 4824 12908 4858
rect 12942 4824 12981 4858
rect 13015 4824 13054 4858
rect 13088 4824 13127 4858
rect 13161 4824 13200 4858
rect 13234 4824 13273 4858
rect 13307 4824 13346 4858
rect -17 4787 17 4824
rect -17 4719 17 4752
rect -17 4651 17 4680
rect -17 4583 17 4608
rect 12564 4758 12598 4824
rect 12564 4690 12598 4724
rect 12564 4622 12598 4656
rect -17 4515 17 4536
rect -17 4447 17 4464
rect 321 4543 345 4581
rect 787 4543 811 4581
rect 321 4437 333 4543
rect 799 4437 811 4543
rect 321 4411 345 4437
rect 787 4411 811 4437
rect 12564 4554 12598 4588
rect 12564 4486 12598 4520
rect 12564 4418 12598 4452
rect -17 4379 17 4392
rect -17 4311 17 4320
rect -17 4243 17 4248
rect -17 4175 17 4176
rect -17 4138 17 4141
rect -17 4066 17 4073
rect -17 3994 17 4005
rect -17 3922 17 3937
rect -17 3850 17 3869
rect 12564 4350 12598 4384
rect 12564 4282 12598 4316
rect 12564 4214 12598 4248
rect 12564 4146 12598 4180
rect 12564 4078 12598 4112
rect 12564 4010 12598 4044
rect 12564 3942 12598 3976
rect 12564 3874 12598 3908
rect -17 3778 17 3801
rect -17 3706 17 3733
rect -17 3634 17 3665
rect 7122 3635 7138 3669
rect 7172 3635 7210 3669
rect 7244 3635 7256 3669
rect 9440 3642 9454 3669
rect 7122 3605 7256 3635
rect 9434 3635 9454 3642
rect 9488 3635 9526 3669
rect 9560 3635 9598 3669
rect 9632 3635 9670 3669
rect 10198 3655 10234 3825
rect 12564 3806 12598 3840
rect 12564 3738 12598 3772
rect 12564 3670 12598 3704
rect -17 3563 17 3597
rect 7538 3561 7552 3567
rect 7586 3561 7624 3595
rect 7885 3580 7896 3595
rect 7658 3561 7672 3567
rect 7930 3561 7968 3595
rect 8002 3580 8019 3595
rect 9132 3580 9144 3595
rect 9178 3561 9216 3595
rect 9250 3580 9266 3595
rect 9434 3582 9704 3635
rect 12564 3602 12598 3636
rect -17 3495 17 3528
rect 8183 3521 8385 3556
rect 10031 3549 10069 3583
rect 10103 3549 10141 3583
rect 8183 3487 8259 3521
rect 8293 3487 8331 3521
rect 8365 3487 8385 3521
rect 8648 3519 8765 3548
rect 8693 3485 8731 3519
rect 12564 3534 12598 3568
rect -17 3427 17 3456
rect -17 3359 17 3393
rect -17 3291 17 3325
rect -17 3223 17 3257
rect -17 3155 17 3189
rect -69 3108 17 3121
rect -35 3087 17 3108
rect 9171 3475 9281 3499
rect 9171 3441 9175 3475
rect 9209 3441 9243 3475
rect 9277 3441 9281 3475
rect 9171 3401 9281 3441
rect 9171 3372 9175 3401
rect 9209 3372 9243 3401
rect 9277 3372 9281 3401
rect 9171 3194 9173 3372
rect 9279 3194 9281 3372
rect 9171 3179 9281 3194
rect 9171 3145 9175 3179
rect 9209 3145 9243 3179
rect 9277 3145 9281 3179
rect 9171 3105 9281 3145
rect -69 3036 -35 3074
rect -69 2964 -35 2992
rect -69 2890 -35 2924
rect 9171 3071 9175 3105
rect 9209 3071 9243 3105
rect 9277 3071 9281 3105
rect 9171 3031 9281 3071
rect 9171 2997 9175 3031
rect 9209 2997 9243 3031
rect 9277 2997 9281 3031
rect 9171 2957 9281 2997
rect 9171 2923 9175 2957
rect 9209 2923 9243 2957
rect 9277 2923 9281 2957
rect 9171 2899 9281 2923
rect 12564 3466 12598 3500
rect 12564 3398 12598 3432
rect 12564 3330 12598 3364
rect 12564 3262 12598 3296
rect 12564 3194 12598 3228
rect 12564 3126 12598 3160
rect 12564 3058 12598 3092
rect 12564 2990 12598 3024
rect 12564 2922 12598 2956
rect -69 2822 -35 2856
rect -69 2754 -35 2788
rect 12564 2854 12598 2888
rect 12564 2786 12598 2820
rect -69 2707 -35 2720
rect -69 2635 -35 2652
rect -69 2563 -35 2584
rect -69 2491 -35 2516
rect -69 2419 -35 2448
rect -69 2347 -35 2380
rect 12564 2718 12598 2752
rect 12564 2650 12598 2684
rect 12564 2582 12598 2616
rect 12564 2514 12598 2548
rect 12564 2446 12598 2480
rect 12564 2378 12598 2412
rect 1095 2341 1134 2375
rect 1168 2341 1207 2375
rect 1241 2341 1280 2375
rect 1314 2341 1353 2375
rect 1387 2341 1426 2375
rect 1460 2341 1499 2375
rect 1533 2341 1572 2375
rect 1606 2341 1645 2375
rect 1679 2341 1718 2375
rect 1752 2341 1791 2375
rect 1825 2341 1864 2375
rect 1898 2341 1937 2375
rect 1971 2341 2010 2375
rect 2044 2341 2083 2375
rect 2117 2341 2156 2375
rect 2190 2341 2229 2375
rect 2263 2341 2302 2375
rect 2336 2341 2375 2375
rect 2409 2341 2448 2375
rect 2482 2341 2521 2375
rect 2555 2341 2594 2375
rect 2628 2341 2667 2375
rect 2701 2341 2740 2375
rect 2774 2341 2813 2375
rect 2847 2341 2886 2375
rect 2920 2341 2959 2375
rect 2993 2341 3032 2375
rect 3066 2341 3105 2375
rect 3139 2341 3178 2375
rect 3212 2341 3251 2375
rect 3285 2341 3324 2375
rect 3358 2341 3397 2375
rect 3431 2341 3470 2375
rect 3504 2341 3543 2375
rect 3577 2341 3616 2375
rect 3650 2341 3689 2375
rect 3723 2341 3762 2375
rect 3796 2341 3835 2375
rect 3869 2341 3907 2375
rect 3941 2341 3979 2375
rect 4013 2341 4051 2375
rect 4085 2341 4123 2375
rect 4157 2341 4195 2375
rect 4229 2341 4267 2375
rect 4301 2341 4339 2375
rect -69 2278 -35 2312
rect 12564 2310 12598 2344
rect -69 2210 -35 2244
rect 10154 2245 10229 2269
rect 10188 2211 10229 2245
rect -69 2142 -35 2176
rect 3176 2174 4464 2182
rect 3176 2140 3200 2174
rect 3234 2140 3271 2174
rect 3305 2140 3342 2174
rect 3376 2140 3413 2174
rect 3447 2140 3484 2174
rect 3518 2140 3555 2174
rect 3589 2140 3626 2174
rect 3660 2140 3697 2174
rect 3731 2140 3768 2174
rect 3802 2140 3839 2174
rect 3873 2140 3910 2174
rect 3944 2140 3981 2174
rect 4015 2140 4052 2174
rect 4086 2140 4123 2174
rect 4157 2140 4194 2174
rect 4228 2140 4265 2174
rect 4299 2140 4336 2174
rect 4370 2140 4406 2174
rect 4440 2140 4464 2174
rect 3176 2132 4464 2140
rect 10154 2177 10229 2211
rect 10188 2143 10229 2177
rect -69 2074 -35 2108
rect -69 2006 -35 2040
rect 3316 2008 3350 2132
rect 3628 2008 3662 2132
rect -69 1938 -35 1972
rect -69 1870 -35 1904
rect -69 1802 -35 1836
rect -69 1734 -35 1768
rect -69 1666 -35 1700
rect -69 1598 -35 1632
rect -69 1530 -35 1564
rect -69 1462 -35 1496
rect -69 1394 -35 1428
rect -69 1326 -35 1360
rect -69 1258 -35 1292
rect -35 1224 661 1244
rect -69 1220 661 1224
rect -69 1190 83 1220
rect -35 1186 83 1190
rect 117 1186 151 1220
rect 185 1186 219 1220
rect 253 1186 287 1220
rect 321 1186 355 1220
rect 389 1186 423 1220
rect 457 1186 491 1220
rect 525 1186 559 1220
rect 593 1186 627 1220
rect -35 1179 661 1186
rect -35 1156 66 1179
rect -69 1145 66 1156
rect 100 1151 141 1179
rect 175 1151 216 1179
rect 250 1151 291 1179
rect 325 1151 367 1179
rect 401 1151 443 1179
rect 477 1151 519 1179
rect 553 1151 595 1179
rect 629 1151 661 1179
rect 117 1145 141 1151
rect 185 1145 216 1151
rect -69 1122 83 1145
rect -35 1117 83 1122
rect 117 1117 151 1145
rect 185 1117 219 1145
rect 253 1117 287 1151
rect 325 1145 355 1151
rect 401 1145 423 1151
rect 477 1145 491 1151
rect 553 1145 559 1151
rect 321 1117 355 1145
rect 389 1117 423 1145
rect 457 1117 491 1145
rect 525 1117 559 1145
rect 593 1145 595 1151
rect 593 1117 627 1145
rect -35 1107 661 1117
rect -35 1088 66 1107
rect -69 1073 66 1088
rect 100 1082 141 1107
rect 175 1082 216 1107
rect 250 1082 291 1107
rect 325 1082 367 1107
rect 401 1082 443 1107
rect 477 1082 519 1107
rect 553 1082 595 1107
rect 629 1082 661 1107
rect 117 1073 141 1082
rect 185 1073 216 1082
rect -69 1054 83 1073
rect -35 1048 83 1054
rect 117 1048 151 1073
rect 185 1048 219 1073
rect 253 1048 287 1082
rect 325 1073 355 1082
rect 401 1073 423 1082
rect 477 1073 491 1082
rect 553 1073 559 1082
rect 321 1048 355 1073
rect 389 1048 423 1073
rect 457 1048 491 1073
rect 525 1048 559 1073
rect 593 1073 595 1082
rect 593 1048 627 1073
rect -35 1035 661 1048
rect -35 1020 66 1035
rect -69 1001 66 1020
rect 100 1013 141 1035
rect 175 1013 216 1035
rect 250 1013 291 1035
rect 325 1013 367 1035
rect 401 1013 443 1035
rect 477 1013 519 1035
rect 553 1013 595 1035
rect 629 1013 661 1035
rect 3940 1008 4072 2132
rect 10154 2109 10229 2143
rect 10188 2075 10229 2109
rect 10154 2041 10229 2075
rect 10188 2007 10229 2041
rect 10154 1973 10229 2007
rect 8463 1930 8701 1954
rect 8497 1896 8531 1930
rect 8565 1896 8599 1930
rect 8633 1896 8667 1930
rect 8463 1856 8701 1896
rect 8497 1822 8531 1856
rect 8565 1822 8599 1856
rect 8633 1822 8667 1856
rect 8463 1782 8701 1822
rect 8497 1748 8531 1782
rect 8565 1748 8599 1782
rect 8633 1748 8667 1782
rect 8463 1708 8701 1748
rect 8497 1674 8531 1708
rect 8565 1674 8599 1708
rect 8633 1674 8667 1708
rect 8463 1634 8701 1674
rect 9155 1930 9221 1954
rect 9155 1896 9171 1930
rect 9205 1896 9221 1930
rect 9155 1829 9221 1896
rect 9155 1795 9171 1829
rect 9205 1795 9221 1829
rect 9155 1728 9221 1795
rect 10188 1939 10229 1973
rect 10154 1905 10229 1939
rect 10188 1871 10229 1905
rect 10154 1837 10229 1871
rect 10188 1803 10229 1837
rect 10154 1779 10229 1803
rect 9155 1723 9171 1728
rect 9205 1723 9221 1728
rect 9205 1694 9227 1723
rect 9189 1689 9227 1694
rect 9155 1670 9221 1689
rect 8497 1600 8531 1634
rect 8565 1600 8599 1634
rect 8633 1600 8667 1634
rect 8463 1560 8701 1600
rect 10195 1564 10229 1779
rect 12564 2242 12598 2276
rect 12564 2174 12598 2208
rect 12564 2106 12598 2140
rect 12564 2038 12598 2072
rect 12564 1970 12598 2004
rect 12564 1902 12598 1936
rect 12564 1834 12598 1868
rect 12564 1766 12598 1800
rect 12591 1708 12598 1732
rect 12557 1698 12598 1708
rect 12557 1670 12564 1698
rect 12591 1636 12598 1664
rect 12557 1630 12598 1636
rect 12557 1598 12564 1630
rect 12591 1564 12598 1596
rect 8497 1526 8531 1560
rect 8565 1526 8599 1560
rect 8633 1526 8667 1560
rect 8463 1487 8701 1526
rect 8497 1453 8531 1487
rect 8565 1453 8599 1487
rect 8633 1453 8667 1487
rect 12564 1562 12598 1564
rect 12564 1494 12598 1528
rect 8463 1414 8701 1453
rect 8497 1380 8531 1414
rect 8565 1380 8599 1414
rect 8633 1380 8667 1414
rect 8463 1341 8701 1380
rect 8497 1307 8531 1341
rect 8565 1307 8599 1341
rect 8633 1307 8667 1341
rect 8463 1268 8701 1307
rect 12591 1440 12598 1460
rect 12557 1426 12598 1440
rect 12557 1402 12564 1426
rect 12591 1368 12598 1392
rect 12557 1358 12598 1368
rect 12557 1330 12564 1358
rect 12591 1296 12598 1324
rect 8497 1234 8531 1268
rect 8565 1234 8599 1268
rect 8633 1234 8667 1268
rect 8463 1221 8701 1234
rect 12564 1290 12598 1296
rect 12564 1222 12598 1256
rect 12564 1154 12598 1188
rect 12564 1086 12598 1120
rect 12564 1018 12598 1052
rect -69 986 83 1001
rect -35 963 83 986
rect -35 952 66 963
rect -69 929 66 952
rect -69 918 83 929
rect -35 891 83 918
rect -35 884 66 891
rect -69 857 66 884
rect -69 850 83 857
rect -35 843 83 850
rect 12564 950 12598 984
rect 12846 932 12932 2350
rect 13000 932 13086 2350
rect 13144 932 13230 2350
rect 12564 898 12598 916
rect 12564 846 12598 848
rect -35 816 661 843
rect -69 814 661 816
rect 12157 826 12598 846
rect 12157 814 12564 826
rect -69 813 12564 814
rect -69 782 12190 813
rect -35 781 12190 782
rect -35 748 121 781
rect -69 747 121 748
rect 155 747 189 781
rect 227 747 257 781
rect 299 747 325 781
rect 371 747 393 781
rect 443 747 461 781
rect 515 747 529 781
rect 587 747 597 781
rect 659 747 665 781
rect 731 747 733 781
rect 767 747 769 781
rect 835 747 841 781
rect 903 747 913 781
rect 971 747 985 781
rect 1039 747 1057 781
rect 1107 747 1129 781
rect 1175 747 1201 781
rect 1243 747 1273 781
rect 1311 747 1345 781
rect 1379 747 1413 781
rect 1451 747 1481 781
rect 1523 747 1549 781
rect 1595 747 1617 781
rect 1667 747 1685 781
rect 1739 747 1753 781
rect 1811 747 1821 781
rect 1883 747 1889 781
rect 1955 747 1957 781
rect 1991 747 1993 781
rect 2059 747 2065 781
rect 2127 747 2137 781
rect 2195 747 2209 781
rect 2263 747 2281 781
rect 2331 747 2353 781
rect 2399 747 2425 781
rect 2467 747 2497 781
rect 2535 747 2569 781
rect 2603 747 2637 781
rect 2675 747 2705 781
rect 2747 747 2773 781
rect 2819 747 2841 781
rect 2891 747 2909 781
rect 2963 747 2977 781
rect 3035 747 3045 781
rect 3107 747 3113 781
rect 3179 747 3181 781
rect 3215 747 3217 781
rect 3283 747 3289 781
rect 3351 747 3361 781
rect 3419 747 3433 781
rect 3487 747 3505 781
rect 3555 747 3577 781
rect 3623 747 3649 781
rect 3691 747 3721 781
rect 3759 747 3793 781
rect 3827 747 3861 781
rect 3899 747 3929 781
rect 3971 747 3997 781
rect 4043 747 4065 781
rect 4115 747 4133 781
rect 4187 747 4201 781
rect 4259 747 4269 781
rect 4331 747 4337 781
rect 4403 747 4405 781
rect 4439 747 4441 781
rect 4507 747 4513 781
rect 4575 747 4585 781
rect 4643 747 4657 781
rect 4711 747 4729 781
rect 4779 747 4801 781
rect 4847 747 4873 781
rect 4915 747 4945 781
rect 4983 747 5017 781
rect 5051 747 5085 781
rect 5123 747 5153 781
rect 5195 747 5221 781
rect 5267 747 5289 781
rect 5339 747 5357 781
rect 5411 747 5425 781
rect 5483 747 5493 781
rect 5555 747 5561 781
rect 5627 747 5629 781
rect 5663 747 5665 781
rect 5731 747 5737 781
rect 5799 747 5809 781
rect 5867 747 5881 781
rect 5935 747 5953 781
rect 6003 747 6025 781
rect 6071 747 6097 781
rect 6139 747 6169 781
rect 6207 747 6241 781
rect 6275 747 6309 781
rect 6347 747 6377 781
rect 6419 747 6445 781
rect 6491 747 6513 781
rect 6563 747 6581 781
rect 6635 747 6649 781
rect 6707 747 6717 781
rect 6779 747 6785 781
rect 6851 747 6853 781
rect 6887 747 6889 781
rect 6955 747 6961 781
rect 7023 747 7033 781
rect 7091 747 7105 781
rect 7159 747 7177 781
rect 7227 747 7249 781
rect 7295 747 7321 781
rect 7363 747 7393 781
rect 7431 747 7465 781
rect 7499 747 7533 781
rect 7571 747 7601 781
rect 7643 747 7669 781
rect 7715 747 7737 781
rect 7787 747 7805 781
rect 7859 747 7873 781
rect 7931 747 7941 781
rect 8003 747 8009 781
rect 8075 747 8077 781
rect 8111 747 8113 781
rect 8179 747 8185 781
rect 8247 747 8257 781
rect 8315 747 8329 781
rect 8383 747 8401 781
rect 8451 747 8473 781
rect 8519 747 8545 781
rect 8587 747 8617 781
rect 8655 747 8689 781
rect 8723 747 8757 781
rect 8795 747 8825 781
rect 8867 747 8893 781
rect 8939 747 8961 781
rect 9011 747 9029 781
rect 9083 747 9097 781
rect 9155 747 9165 781
rect 9227 747 9233 781
rect 9299 747 9301 781
rect 9335 747 9337 781
rect 9403 747 9409 781
rect 9471 747 9481 781
rect 9539 747 9553 781
rect 9607 747 9625 781
rect 9675 747 9697 781
rect 9743 747 9769 781
rect 9811 747 9841 781
rect 9879 747 9913 781
rect 9947 747 9981 781
rect 10019 747 10049 781
rect 10091 747 10117 781
rect 10163 747 10185 781
rect 10235 747 10253 781
rect 10307 747 10321 781
rect 10379 747 10389 781
rect 10451 747 10457 781
rect 10523 747 10525 781
rect 10559 747 10561 781
rect 10627 747 10633 781
rect 10695 747 10705 781
rect 10763 747 10777 781
rect 10831 747 10849 781
rect 10899 747 10921 781
rect 10967 747 10993 781
rect 11035 747 11065 781
rect 11103 747 11137 781
rect 11171 747 11205 781
rect 11243 747 11273 781
rect 11315 747 11341 781
rect 11387 747 11409 781
rect 11459 747 11477 781
rect 11531 747 11545 781
rect 11603 747 11613 781
rect 11675 747 11681 781
rect 11747 747 11749 781
rect 11783 747 11785 781
rect 11851 747 11857 781
rect 11919 747 11929 781
rect 11987 747 12001 781
rect 12055 747 12073 781
rect 12123 779 12190 781
rect 12224 779 12258 813
rect 12296 779 12326 813
rect 12368 779 12394 813
rect 12440 779 12462 813
rect 12512 780 12564 813
rect 12512 779 12598 780
rect 12123 747 12598 779
rect -69 746 12598 747
rect -69 714 12257 746
<< viali >>
rect -17 4824 17 4858
rect 55 4824 89 4858
rect 127 4824 161 4858
rect 199 4824 229 4858
rect 229 4824 233 4858
rect 271 4824 297 4858
rect 297 4824 305 4858
rect 343 4824 365 4858
rect 365 4824 377 4858
rect 415 4824 433 4858
rect 433 4824 449 4858
rect 508 4824 535 4858
rect 535 4824 542 4858
rect 580 4824 603 4858
rect 603 4824 614 4858
rect 652 4824 671 4858
rect 671 4824 686 4858
rect 724 4824 739 4858
rect 739 4824 758 4858
rect 796 4824 807 4858
rect 807 4824 830 4858
rect 868 4824 875 4858
rect 875 4824 902 4858
rect 940 4824 943 4858
rect 943 4824 974 4858
rect 1012 4824 1045 4858
rect 1045 4824 1046 4858
rect 1084 4824 1113 4858
rect 1113 4824 1118 4858
rect 1156 4824 1181 4858
rect 1181 4824 1190 4858
rect 1228 4824 1249 4858
rect 1249 4824 1262 4858
rect 1300 4824 1317 4858
rect 1317 4824 1334 4858
rect 1372 4824 1385 4858
rect 1385 4824 1406 4858
rect 1444 4824 1453 4858
rect 1453 4824 1478 4858
rect 1516 4824 1521 4858
rect 1521 4824 1550 4858
rect 1588 4824 1589 4858
rect 1589 4824 1622 4858
rect 1660 4824 1691 4858
rect 1691 4824 1694 4858
rect 1732 4824 1759 4858
rect 1759 4824 1766 4858
rect 1804 4824 1827 4858
rect 1827 4824 1838 4858
rect 1876 4824 1895 4858
rect 1895 4824 1910 4858
rect 1948 4824 1963 4858
rect 1963 4824 1982 4858
rect 2020 4824 2031 4858
rect 2031 4824 2054 4858
rect 2092 4824 2099 4858
rect 2099 4824 2126 4858
rect 2164 4824 2167 4858
rect 2167 4824 2198 4858
rect 2236 4824 2269 4858
rect 2269 4824 2270 4858
rect 2308 4824 2337 4858
rect 2337 4824 2342 4858
rect 2380 4824 2405 4858
rect 2405 4824 2414 4858
rect 2452 4824 2473 4858
rect 2473 4824 2486 4858
rect 2524 4824 2541 4858
rect 2541 4824 2558 4858
rect 2596 4824 2609 4858
rect 2609 4824 2630 4858
rect 2668 4824 2677 4858
rect 2677 4824 2702 4858
rect 2740 4824 2745 4858
rect 2745 4824 2774 4858
rect 2812 4824 2813 4858
rect 2813 4824 2846 4858
rect 2884 4824 2915 4858
rect 2915 4824 2918 4858
rect 2956 4824 2983 4858
rect 2983 4824 2990 4858
rect 3028 4824 3051 4858
rect 3051 4824 3062 4858
rect 3100 4824 3119 4858
rect 3119 4824 3134 4858
rect 3172 4824 3187 4858
rect 3187 4824 3206 4858
rect 3244 4824 3255 4858
rect 3255 4824 3278 4858
rect 3316 4824 3323 4858
rect 3323 4824 3350 4858
rect 3388 4824 3391 4858
rect 3391 4824 3422 4858
rect 3460 4824 3493 4858
rect 3493 4824 3494 4858
rect 3532 4824 3561 4858
rect 3561 4824 3566 4858
rect 3604 4824 3629 4858
rect 3629 4824 3638 4858
rect 3676 4824 3697 4858
rect 3697 4824 3710 4858
rect 3748 4824 3765 4858
rect 3765 4824 3782 4858
rect 3820 4824 3833 4858
rect 3833 4824 3854 4858
rect 3892 4824 3901 4858
rect 3901 4824 3926 4858
rect 3964 4824 3969 4858
rect 3969 4824 3998 4858
rect 4036 4824 4037 4858
rect 4037 4824 4070 4858
rect 4108 4824 4139 4858
rect 4139 4824 4142 4858
rect 4180 4824 4207 4858
rect 4207 4824 4214 4858
rect 4252 4824 4275 4858
rect 4275 4824 4286 4858
rect 4324 4824 4343 4858
rect 4343 4824 4358 4858
rect 4396 4824 4411 4858
rect 4411 4824 4430 4858
rect 4468 4824 4479 4858
rect 4479 4824 4502 4858
rect 4540 4824 4547 4858
rect 4547 4824 4574 4858
rect 4612 4824 4615 4858
rect 4615 4824 4646 4858
rect 4684 4824 4717 4858
rect 4717 4824 4718 4858
rect 4756 4824 4785 4858
rect 4785 4824 4790 4858
rect 4828 4824 4853 4858
rect 4853 4824 4862 4858
rect 4900 4824 4921 4858
rect 4921 4824 4934 4858
rect 4972 4824 4989 4858
rect 4989 4824 5006 4858
rect 5044 4824 5057 4858
rect 5057 4824 5078 4858
rect 5116 4824 5125 4858
rect 5125 4824 5150 4858
rect 5188 4824 5193 4858
rect 5193 4824 5222 4858
rect 5260 4824 5261 4858
rect 5261 4824 5294 4858
rect 5332 4824 5363 4858
rect 5363 4824 5366 4858
rect 5404 4824 5431 4858
rect 5431 4824 5438 4858
rect 5476 4824 5499 4858
rect 5499 4824 5510 4858
rect 5548 4824 5567 4858
rect 5567 4824 5582 4858
rect 5620 4824 5635 4858
rect 5635 4824 5654 4858
rect 5692 4824 5703 4858
rect 5703 4824 5726 4858
rect 5764 4824 5771 4858
rect 5771 4824 5798 4858
rect 5836 4824 5839 4858
rect 5839 4824 5870 4858
rect 5908 4824 5941 4858
rect 5941 4824 5942 4858
rect 5980 4824 6009 4858
rect 6009 4824 6014 4858
rect 6052 4824 6077 4858
rect 6077 4824 6086 4858
rect 6124 4824 6145 4858
rect 6145 4824 6158 4858
rect 6196 4824 6213 4858
rect 6213 4824 6230 4858
rect 6268 4824 6281 4858
rect 6281 4824 6302 4858
rect 6340 4824 6349 4858
rect 6349 4824 6374 4858
rect 6412 4824 6417 4858
rect 6417 4824 6446 4858
rect 6484 4824 6485 4858
rect 6485 4824 6518 4858
rect 6556 4824 6587 4858
rect 6587 4824 6590 4858
rect 6628 4824 6655 4858
rect 6655 4824 6662 4858
rect 6700 4824 6723 4858
rect 6723 4824 6734 4858
rect 6772 4824 6791 4858
rect 6791 4824 6806 4858
rect 6844 4824 6859 4858
rect 6859 4824 6878 4858
rect 6916 4824 6927 4858
rect 6927 4824 6950 4858
rect 6988 4824 6995 4858
rect 6995 4824 7022 4858
rect 7060 4824 7063 4858
rect 7063 4824 7094 4858
rect 7132 4824 7165 4858
rect 7165 4824 7166 4858
rect 7204 4824 7233 4858
rect 7233 4824 7238 4858
rect 7276 4824 7301 4858
rect 7301 4824 7310 4858
rect 7348 4824 7369 4858
rect 7369 4824 7382 4858
rect 7420 4824 7437 4858
rect 7437 4824 7454 4858
rect 7492 4824 7505 4858
rect 7505 4824 7526 4858
rect 7564 4824 7573 4858
rect 7573 4824 7598 4858
rect 7636 4824 7641 4858
rect 7641 4824 7670 4858
rect 7708 4824 7709 4858
rect 7709 4824 7742 4858
rect 7780 4824 7811 4858
rect 7811 4824 7814 4858
rect 7852 4824 7879 4858
rect 7879 4824 7886 4858
rect 7924 4824 7947 4858
rect 7947 4824 7958 4858
rect 7996 4824 8015 4858
rect 8015 4824 8030 4858
rect 8068 4824 8083 4858
rect 8083 4824 8102 4858
rect 8140 4824 8151 4858
rect 8151 4824 8174 4858
rect 8212 4824 8219 4858
rect 8219 4824 8246 4858
rect 8284 4824 8287 4858
rect 8287 4824 8318 4858
rect 8356 4824 8389 4858
rect 8389 4824 8390 4858
rect 8428 4824 8457 4858
rect 8457 4824 8462 4858
rect 8500 4824 8525 4858
rect 8525 4824 8534 4858
rect 8572 4824 8593 4858
rect 8593 4824 8606 4858
rect 8644 4824 8661 4858
rect 8661 4824 8678 4858
rect 8716 4824 8729 4858
rect 8729 4824 8750 4858
rect 8788 4824 8797 4858
rect 8797 4824 8822 4858
rect 8860 4824 8865 4858
rect 8865 4824 8894 4858
rect 8932 4824 8933 4858
rect 8933 4824 8966 4858
rect 9004 4824 9035 4858
rect 9035 4824 9038 4858
rect 9076 4824 9103 4858
rect 9103 4824 9110 4858
rect 9148 4824 9171 4858
rect 9171 4824 9182 4858
rect 9220 4824 9239 4858
rect 9239 4824 9254 4858
rect 9292 4824 9307 4858
rect 9307 4824 9326 4858
rect 9364 4824 9375 4858
rect 9375 4824 9398 4858
rect 9436 4824 9443 4858
rect 9443 4824 9470 4858
rect 9508 4824 9511 4858
rect 9511 4824 9542 4858
rect 9580 4824 9613 4858
rect 9613 4824 9614 4858
rect 9652 4824 9681 4858
rect 9681 4824 9686 4858
rect 9724 4824 9749 4858
rect 9749 4824 9758 4858
rect 9796 4824 9817 4858
rect 9817 4824 9830 4858
rect 9868 4824 9885 4858
rect 9885 4824 9902 4858
rect 9940 4824 9953 4858
rect 9953 4824 9974 4858
rect 10012 4824 10021 4858
rect 10021 4824 10046 4858
rect 10084 4824 10089 4858
rect 10089 4824 10118 4858
rect 10156 4824 10157 4858
rect 10157 4824 10190 4858
rect 10228 4824 10259 4858
rect 10259 4824 10262 4858
rect 10300 4824 10327 4858
rect 10327 4824 10334 4858
rect 10372 4824 10395 4858
rect 10395 4824 10406 4858
rect 10444 4824 10463 4858
rect 10463 4824 10478 4858
rect 10516 4824 10531 4858
rect 10531 4824 10550 4858
rect 10588 4824 10599 4858
rect 10599 4824 10622 4858
rect 10660 4824 10667 4858
rect 10667 4824 10694 4858
rect 10732 4824 10735 4858
rect 10735 4824 10766 4858
rect 10804 4824 10837 4858
rect 10837 4824 10838 4858
rect 10876 4824 10905 4858
rect 10905 4824 10910 4858
rect 10948 4824 10973 4858
rect 10973 4824 10982 4858
rect 11020 4824 11041 4858
rect 11041 4824 11054 4858
rect 11092 4824 11109 4858
rect 11109 4824 11126 4858
rect 11164 4824 11177 4858
rect 11177 4824 11198 4858
rect 11236 4824 11245 4858
rect 11245 4824 11270 4858
rect 11308 4824 11313 4858
rect 11313 4824 11342 4858
rect 11380 4824 11381 4858
rect 11381 4824 11414 4858
rect 11452 4824 11483 4858
rect 11483 4824 11486 4858
rect 11524 4824 11551 4858
rect 11551 4824 11558 4858
rect 11596 4824 11619 4858
rect 11619 4824 11630 4858
rect 11668 4824 11687 4858
rect 11687 4824 11702 4858
rect 11740 4824 11755 4858
rect 11755 4824 11774 4858
rect 11813 4824 11823 4858
rect 11823 4824 11847 4858
rect 11886 4824 11891 4858
rect 11891 4824 11920 4858
rect 11959 4824 11993 4858
rect 12032 4824 12061 4858
rect 12061 4824 12066 4858
rect 12105 4824 12129 4858
rect 12129 4824 12139 4858
rect 12178 4824 12197 4858
rect 12197 4824 12212 4858
rect 12251 4824 12265 4858
rect 12265 4824 12285 4858
rect 12324 4824 12333 4858
rect 12333 4824 12358 4858
rect 12397 4824 12401 4858
rect 12401 4824 12431 4858
rect 12470 4824 12504 4858
rect 12543 4824 12577 4858
rect 12616 4824 12650 4858
rect 12689 4824 12723 4858
rect 12762 4824 12796 4858
rect 12835 4824 12869 4858
rect 12908 4824 12942 4858
rect 12981 4824 13015 4858
rect 13054 4824 13088 4858
rect 13127 4824 13161 4858
rect 13200 4824 13234 4858
rect 13273 4824 13307 4858
rect 13346 4824 13380 4858
rect -17 4753 17 4786
rect -17 4752 17 4753
rect -17 4685 17 4714
rect -17 4680 17 4685
rect -17 4617 17 4642
rect -17 4608 17 4617
rect -17 4549 17 4570
rect -17 4536 17 4549
rect -17 4481 17 4498
rect -17 4464 17 4481
rect -17 4413 17 4426
rect -17 4392 17 4413
rect 333 4437 345 4543
rect 345 4437 787 4543
rect 787 4437 799 4543
rect -17 4345 17 4354
rect -17 4320 17 4345
rect -17 4277 17 4282
rect -17 4248 17 4277
rect -17 4209 17 4210
rect -17 4176 17 4209
rect -17 4107 17 4138
rect -17 4104 17 4107
rect -17 4039 17 4066
rect -17 4032 17 4039
rect -17 3971 17 3994
rect -17 3960 17 3971
rect -17 3903 17 3922
rect -17 3888 17 3903
rect -17 3835 17 3850
rect -17 3816 17 3835
rect -17 3767 17 3778
rect -17 3744 17 3767
rect -17 3699 17 3706
rect -17 3672 17 3699
rect -17 3631 17 3634
rect -17 3600 17 3631
rect 7138 3635 7172 3669
rect 7210 3635 7244 3669
rect 9454 3635 9488 3669
rect 9526 3635 9560 3669
rect 9598 3635 9632 3669
rect 9670 3635 9704 3669
rect -17 3529 17 3562
rect 7552 3561 7586 3595
rect 7624 3561 7658 3595
rect 7896 3561 7930 3595
rect 7968 3561 8002 3595
rect 9144 3561 9178 3595
rect 9216 3561 9250 3595
rect -17 3528 17 3529
rect -17 3461 17 3490
rect 9997 3549 10031 3583
rect 10069 3549 10103 3583
rect 10141 3549 10175 3583
rect 8259 3487 8293 3521
rect 8331 3487 8365 3521
rect 8659 3485 8693 3519
rect 8731 3485 8765 3519
rect -17 3456 17 3461
rect -69 3074 -35 3108
rect 9173 3367 9175 3372
rect 9175 3367 9209 3372
rect 9209 3367 9243 3372
rect 9243 3367 9277 3372
rect 9277 3367 9279 3372
rect 9173 3327 9279 3367
rect 9173 3293 9175 3327
rect 9175 3293 9209 3327
rect 9209 3293 9243 3327
rect 9243 3293 9277 3327
rect 9277 3293 9279 3327
rect 9173 3253 9279 3293
rect 9173 3219 9175 3253
rect 9175 3219 9209 3253
rect 9209 3219 9243 3253
rect 9243 3219 9277 3253
rect 9277 3219 9279 3253
rect 9173 3194 9279 3219
rect -69 3026 -35 3036
rect -69 3002 -35 3026
rect -69 2958 -35 2964
rect -69 2930 -35 2958
rect 400 2777 1010 2883
rect -69 2686 -35 2707
rect -69 2673 -35 2686
rect -69 2618 -35 2635
rect -69 2601 -35 2618
rect -69 2550 -35 2563
rect -69 2529 -35 2550
rect -69 2482 -35 2491
rect -69 2457 -35 2482
rect -69 2414 -35 2419
rect -69 2385 -35 2414
rect -69 2346 -35 2347
rect -69 2313 -35 2346
rect 1061 2341 1095 2375
rect 1134 2341 1168 2375
rect 1207 2341 1241 2375
rect 1280 2341 1314 2375
rect 1353 2341 1387 2375
rect 1426 2341 1460 2375
rect 1499 2341 1533 2375
rect 1572 2341 1606 2375
rect 1645 2341 1679 2375
rect 1718 2341 1752 2375
rect 1791 2341 1825 2375
rect 1864 2341 1898 2375
rect 1937 2341 1971 2375
rect 2010 2341 2044 2375
rect 2083 2341 2117 2375
rect 2156 2341 2190 2375
rect 2229 2341 2263 2375
rect 2302 2341 2336 2375
rect 2375 2341 2409 2375
rect 2448 2341 2482 2375
rect 2521 2341 2555 2375
rect 2594 2341 2628 2375
rect 2667 2341 2701 2375
rect 2740 2341 2774 2375
rect 2813 2341 2847 2375
rect 2886 2341 2920 2375
rect 2959 2341 2993 2375
rect 3032 2341 3066 2375
rect 3105 2341 3139 2375
rect 3178 2341 3212 2375
rect 3251 2341 3285 2375
rect 3324 2341 3358 2375
rect 3397 2341 3431 2375
rect 3470 2341 3504 2375
rect 3543 2341 3577 2375
rect 3616 2341 3650 2375
rect 3689 2341 3723 2375
rect 3762 2341 3796 2375
rect 3835 2341 3869 2375
rect 3907 2341 3941 2375
rect 3979 2341 4013 2375
rect 4051 2341 4085 2375
rect 4123 2341 4157 2375
rect 4195 2341 4229 2375
rect 4267 2341 4301 2375
rect 4339 2341 4373 2375
rect 66 1151 100 1179
rect 141 1151 175 1179
rect 216 1151 250 1179
rect 291 1151 325 1179
rect 367 1151 401 1179
rect 443 1151 477 1179
rect 519 1151 553 1179
rect 595 1151 629 1179
rect 66 1145 83 1151
rect 83 1145 100 1151
rect 141 1145 151 1151
rect 151 1145 175 1151
rect 216 1145 219 1151
rect 219 1145 250 1151
rect 291 1145 321 1151
rect 321 1145 325 1151
rect 367 1145 389 1151
rect 389 1145 401 1151
rect 443 1145 457 1151
rect 457 1145 477 1151
rect 519 1145 525 1151
rect 525 1145 553 1151
rect 595 1145 627 1151
rect 627 1145 629 1151
rect 66 1082 100 1107
rect 141 1082 175 1107
rect 216 1082 250 1107
rect 291 1082 325 1107
rect 367 1082 401 1107
rect 443 1082 477 1107
rect 519 1082 553 1107
rect 595 1082 629 1107
rect 66 1073 83 1082
rect 83 1073 100 1082
rect 141 1073 151 1082
rect 151 1073 175 1082
rect 216 1073 219 1082
rect 219 1073 250 1082
rect 291 1073 321 1082
rect 321 1073 325 1082
rect 367 1073 389 1082
rect 389 1073 401 1082
rect 443 1073 457 1082
rect 457 1073 477 1082
rect 519 1073 525 1082
rect 525 1073 553 1082
rect 595 1073 627 1082
rect 627 1073 629 1082
rect 66 1013 100 1035
rect 141 1013 175 1035
rect 216 1013 250 1035
rect 291 1013 325 1035
rect 367 1013 401 1035
rect 443 1013 477 1035
rect 519 1013 553 1035
rect 595 1013 629 1035
rect 66 1001 83 1013
rect 83 1001 100 1013
rect 141 1001 175 1013
rect 216 1001 250 1013
rect 291 1001 325 1013
rect 367 1001 401 1013
rect 443 1001 477 1013
rect 519 1001 553 1013
rect 595 1001 629 1013
rect 9155 1694 9171 1723
rect 9171 1694 9189 1723
rect 9155 1689 9189 1694
rect 9227 1689 9261 1723
rect 12557 1732 12564 1742
rect 12564 1732 12591 1742
rect 12557 1708 12591 1732
rect 12557 1664 12564 1670
rect 12564 1664 12591 1670
rect 12557 1636 12591 1664
rect 12557 1596 12564 1598
rect 12564 1596 12591 1598
rect 12557 1564 12591 1596
rect 12557 1460 12564 1474
rect 12564 1460 12591 1474
rect 12557 1440 12591 1460
rect 12557 1392 12564 1402
rect 12564 1392 12591 1402
rect 12557 1368 12591 1392
rect 12557 1324 12564 1330
rect 12564 1324 12591 1330
rect 12557 1296 12591 1324
rect 8463 1195 8713 1221
rect 8463 1161 8497 1195
rect 8497 1161 8531 1195
rect 8531 1161 8565 1195
rect 8565 1161 8599 1195
rect 8599 1161 8633 1195
rect 8633 1161 8667 1195
rect 8667 1161 8701 1195
rect 8701 1161 8713 1195
rect 8463 1122 8713 1161
rect 8463 1088 8497 1122
rect 8497 1088 8531 1122
rect 8531 1088 8565 1122
rect 8565 1088 8599 1122
rect 8599 1088 8633 1122
rect 8633 1088 8667 1122
rect 8667 1088 8701 1122
rect 8701 1088 8713 1122
rect 8463 1043 8713 1088
rect 66 929 83 963
rect 83 929 100 963
rect 141 929 175 963
rect 216 929 250 963
rect 291 929 325 963
rect 367 929 401 963
rect 443 929 477 963
rect 519 929 553 963
rect 595 929 629 963
rect 66 857 83 891
rect 83 857 100 891
rect 141 857 175 891
rect 216 857 250 891
rect 291 857 325 891
rect 367 857 401 891
rect 443 857 477 891
rect 519 857 553 891
rect 595 857 629 891
rect 12564 882 12598 898
rect 12564 864 12598 882
rect 12564 814 12598 826
rect 121 747 155 781
rect 193 747 223 781
rect 223 747 227 781
rect 265 747 291 781
rect 291 747 299 781
rect 337 747 359 781
rect 359 747 371 781
rect 409 747 427 781
rect 427 747 443 781
rect 481 747 495 781
rect 495 747 515 781
rect 553 747 563 781
rect 563 747 587 781
rect 625 747 631 781
rect 631 747 659 781
rect 697 747 699 781
rect 699 747 731 781
rect 769 747 801 781
rect 801 747 803 781
rect 841 747 869 781
rect 869 747 875 781
rect 913 747 937 781
rect 937 747 947 781
rect 985 747 1005 781
rect 1005 747 1019 781
rect 1057 747 1073 781
rect 1073 747 1091 781
rect 1129 747 1141 781
rect 1141 747 1163 781
rect 1201 747 1209 781
rect 1209 747 1235 781
rect 1273 747 1277 781
rect 1277 747 1307 781
rect 1345 747 1379 781
rect 1417 747 1447 781
rect 1447 747 1451 781
rect 1489 747 1515 781
rect 1515 747 1523 781
rect 1561 747 1583 781
rect 1583 747 1595 781
rect 1633 747 1651 781
rect 1651 747 1667 781
rect 1705 747 1719 781
rect 1719 747 1739 781
rect 1777 747 1787 781
rect 1787 747 1811 781
rect 1849 747 1855 781
rect 1855 747 1883 781
rect 1921 747 1923 781
rect 1923 747 1955 781
rect 1993 747 2025 781
rect 2025 747 2027 781
rect 2065 747 2093 781
rect 2093 747 2099 781
rect 2137 747 2161 781
rect 2161 747 2171 781
rect 2209 747 2229 781
rect 2229 747 2243 781
rect 2281 747 2297 781
rect 2297 747 2315 781
rect 2353 747 2365 781
rect 2365 747 2387 781
rect 2425 747 2433 781
rect 2433 747 2459 781
rect 2497 747 2501 781
rect 2501 747 2531 781
rect 2569 747 2603 781
rect 2641 747 2671 781
rect 2671 747 2675 781
rect 2713 747 2739 781
rect 2739 747 2747 781
rect 2785 747 2807 781
rect 2807 747 2819 781
rect 2857 747 2875 781
rect 2875 747 2891 781
rect 2929 747 2943 781
rect 2943 747 2963 781
rect 3001 747 3011 781
rect 3011 747 3035 781
rect 3073 747 3079 781
rect 3079 747 3107 781
rect 3145 747 3147 781
rect 3147 747 3179 781
rect 3217 747 3249 781
rect 3249 747 3251 781
rect 3289 747 3317 781
rect 3317 747 3323 781
rect 3361 747 3385 781
rect 3385 747 3395 781
rect 3433 747 3453 781
rect 3453 747 3467 781
rect 3505 747 3521 781
rect 3521 747 3539 781
rect 3577 747 3589 781
rect 3589 747 3611 781
rect 3649 747 3657 781
rect 3657 747 3683 781
rect 3721 747 3725 781
rect 3725 747 3755 781
rect 3793 747 3827 781
rect 3865 747 3895 781
rect 3895 747 3899 781
rect 3937 747 3963 781
rect 3963 747 3971 781
rect 4009 747 4031 781
rect 4031 747 4043 781
rect 4081 747 4099 781
rect 4099 747 4115 781
rect 4153 747 4167 781
rect 4167 747 4187 781
rect 4225 747 4235 781
rect 4235 747 4259 781
rect 4297 747 4303 781
rect 4303 747 4331 781
rect 4369 747 4371 781
rect 4371 747 4403 781
rect 4441 747 4473 781
rect 4473 747 4475 781
rect 4513 747 4541 781
rect 4541 747 4547 781
rect 4585 747 4609 781
rect 4609 747 4619 781
rect 4657 747 4677 781
rect 4677 747 4691 781
rect 4729 747 4745 781
rect 4745 747 4763 781
rect 4801 747 4813 781
rect 4813 747 4835 781
rect 4873 747 4881 781
rect 4881 747 4907 781
rect 4945 747 4949 781
rect 4949 747 4979 781
rect 5017 747 5051 781
rect 5089 747 5119 781
rect 5119 747 5123 781
rect 5161 747 5187 781
rect 5187 747 5195 781
rect 5233 747 5255 781
rect 5255 747 5267 781
rect 5305 747 5323 781
rect 5323 747 5339 781
rect 5377 747 5391 781
rect 5391 747 5411 781
rect 5449 747 5459 781
rect 5459 747 5483 781
rect 5521 747 5527 781
rect 5527 747 5555 781
rect 5593 747 5595 781
rect 5595 747 5627 781
rect 5665 747 5697 781
rect 5697 747 5699 781
rect 5737 747 5765 781
rect 5765 747 5771 781
rect 5809 747 5833 781
rect 5833 747 5843 781
rect 5881 747 5901 781
rect 5901 747 5915 781
rect 5953 747 5969 781
rect 5969 747 5987 781
rect 6025 747 6037 781
rect 6037 747 6059 781
rect 6097 747 6105 781
rect 6105 747 6131 781
rect 6169 747 6173 781
rect 6173 747 6203 781
rect 6241 747 6275 781
rect 6313 747 6343 781
rect 6343 747 6347 781
rect 6385 747 6411 781
rect 6411 747 6419 781
rect 6457 747 6479 781
rect 6479 747 6491 781
rect 6529 747 6547 781
rect 6547 747 6563 781
rect 6601 747 6615 781
rect 6615 747 6635 781
rect 6673 747 6683 781
rect 6683 747 6707 781
rect 6745 747 6751 781
rect 6751 747 6779 781
rect 6817 747 6819 781
rect 6819 747 6851 781
rect 6889 747 6921 781
rect 6921 747 6923 781
rect 6961 747 6989 781
rect 6989 747 6995 781
rect 7033 747 7057 781
rect 7057 747 7067 781
rect 7105 747 7125 781
rect 7125 747 7139 781
rect 7177 747 7193 781
rect 7193 747 7211 781
rect 7249 747 7261 781
rect 7261 747 7283 781
rect 7321 747 7329 781
rect 7329 747 7355 781
rect 7393 747 7397 781
rect 7397 747 7427 781
rect 7465 747 7499 781
rect 7537 747 7567 781
rect 7567 747 7571 781
rect 7609 747 7635 781
rect 7635 747 7643 781
rect 7681 747 7703 781
rect 7703 747 7715 781
rect 7753 747 7771 781
rect 7771 747 7787 781
rect 7825 747 7839 781
rect 7839 747 7859 781
rect 7897 747 7907 781
rect 7907 747 7931 781
rect 7969 747 7975 781
rect 7975 747 8003 781
rect 8041 747 8043 781
rect 8043 747 8075 781
rect 8113 747 8145 781
rect 8145 747 8147 781
rect 8185 747 8213 781
rect 8213 747 8219 781
rect 8257 747 8281 781
rect 8281 747 8291 781
rect 8329 747 8349 781
rect 8349 747 8363 781
rect 8401 747 8417 781
rect 8417 747 8435 781
rect 8473 747 8485 781
rect 8485 747 8507 781
rect 8545 747 8553 781
rect 8553 747 8579 781
rect 8617 747 8621 781
rect 8621 747 8651 781
rect 8689 747 8723 781
rect 8761 747 8791 781
rect 8791 747 8795 781
rect 8833 747 8859 781
rect 8859 747 8867 781
rect 8905 747 8927 781
rect 8927 747 8939 781
rect 8977 747 8995 781
rect 8995 747 9011 781
rect 9049 747 9063 781
rect 9063 747 9083 781
rect 9121 747 9131 781
rect 9131 747 9155 781
rect 9193 747 9199 781
rect 9199 747 9227 781
rect 9265 747 9267 781
rect 9267 747 9299 781
rect 9337 747 9369 781
rect 9369 747 9371 781
rect 9409 747 9437 781
rect 9437 747 9443 781
rect 9481 747 9505 781
rect 9505 747 9515 781
rect 9553 747 9573 781
rect 9573 747 9587 781
rect 9625 747 9641 781
rect 9641 747 9659 781
rect 9697 747 9709 781
rect 9709 747 9731 781
rect 9769 747 9777 781
rect 9777 747 9803 781
rect 9841 747 9845 781
rect 9845 747 9875 781
rect 9913 747 9947 781
rect 9985 747 10015 781
rect 10015 747 10019 781
rect 10057 747 10083 781
rect 10083 747 10091 781
rect 10129 747 10151 781
rect 10151 747 10163 781
rect 10201 747 10219 781
rect 10219 747 10235 781
rect 10273 747 10287 781
rect 10287 747 10307 781
rect 10345 747 10355 781
rect 10355 747 10379 781
rect 10417 747 10423 781
rect 10423 747 10451 781
rect 10489 747 10491 781
rect 10491 747 10523 781
rect 10561 747 10593 781
rect 10593 747 10595 781
rect 10633 747 10661 781
rect 10661 747 10667 781
rect 10705 747 10729 781
rect 10729 747 10739 781
rect 10777 747 10797 781
rect 10797 747 10811 781
rect 10849 747 10865 781
rect 10865 747 10883 781
rect 10921 747 10933 781
rect 10933 747 10955 781
rect 10993 747 11001 781
rect 11001 747 11027 781
rect 11065 747 11069 781
rect 11069 747 11099 781
rect 11137 747 11171 781
rect 11209 747 11239 781
rect 11239 747 11243 781
rect 11281 747 11307 781
rect 11307 747 11315 781
rect 11353 747 11375 781
rect 11375 747 11387 781
rect 11425 747 11443 781
rect 11443 747 11459 781
rect 11497 747 11511 781
rect 11511 747 11531 781
rect 11569 747 11579 781
rect 11579 747 11603 781
rect 11641 747 11647 781
rect 11647 747 11675 781
rect 11713 747 11715 781
rect 11715 747 11747 781
rect 11785 747 11817 781
rect 11817 747 11819 781
rect 11857 747 11885 781
rect 11885 747 11891 781
rect 11929 747 11953 781
rect 11953 747 11963 781
rect 12001 747 12021 781
rect 12021 747 12035 781
rect 12073 747 12089 781
rect 12089 747 12107 781
rect 12190 779 12224 813
rect 12262 779 12292 813
rect 12292 779 12296 813
rect 12334 779 12360 813
rect 12360 779 12368 813
rect 12406 779 12428 813
rect 12428 779 12440 813
rect 12478 779 12496 813
rect 12496 779 12512 813
rect 12564 792 12598 814
<< metal1 >>
rect -26 4867 32 4870
tri 32 4867 35 4870 sw
rect -26 4864 35 4867
tri 35 4864 38 4867 sw
rect -26 4858 13392 4864
rect -26 4824 -17 4858
rect 17 4824 55 4858
rect 89 4824 127 4858
rect 161 4824 199 4858
rect 233 4824 271 4858
rect 305 4824 343 4858
rect 377 4824 415 4858
rect 449 4824 508 4858
rect 542 4824 580 4858
rect 614 4824 652 4858
rect 686 4824 724 4858
rect 758 4824 796 4858
rect 830 4824 868 4858
rect 902 4824 940 4858
rect 974 4824 1012 4858
rect 1046 4824 1084 4858
rect 1118 4824 1156 4858
rect 1190 4824 1228 4858
rect 1262 4824 1300 4858
rect 1334 4824 1372 4858
rect 1406 4824 1444 4858
rect 1478 4824 1516 4858
rect 1550 4824 1588 4858
rect 1622 4824 1660 4858
rect 1694 4824 1732 4858
rect 1766 4824 1804 4858
rect 1838 4824 1876 4858
rect 1910 4824 1948 4858
rect 1982 4824 2020 4858
rect 2054 4824 2092 4858
rect 2126 4824 2164 4858
rect 2198 4824 2236 4858
rect 2270 4824 2308 4858
rect 2342 4824 2380 4858
rect 2414 4824 2452 4858
rect 2486 4824 2524 4858
rect 2558 4824 2596 4858
rect 2630 4824 2668 4858
rect 2702 4824 2740 4858
rect 2774 4824 2812 4858
rect 2846 4824 2884 4858
rect 2918 4824 2956 4858
rect 2990 4824 3028 4858
rect 3062 4824 3100 4858
rect 3134 4824 3172 4858
rect 3206 4824 3244 4858
rect 3278 4824 3316 4858
rect 3350 4824 3388 4858
rect 3422 4824 3460 4858
rect 3494 4824 3532 4858
rect 3566 4824 3604 4858
rect 3638 4824 3676 4858
rect 3710 4824 3748 4858
rect 3782 4824 3820 4858
rect 3854 4824 3892 4858
rect 3926 4824 3964 4858
rect 3998 4824 4036 4858
rect 4070 4824 4108 4858
rect 4142 4824 4180 4858
rect 4214 4824 4252 4858
rect 4286 4824 4324 4858
rect 4358 4824 4396 4858
rect 4430 4824 4468 4858
rect 4502 4824 4540 4858
rect 4574 4824 4612 4858
rect 4646 4824 4684 4858
rect 4718 4824 4756 4858
rect 4790 4824 4828 4858
rect 4862 4824 4900 4858
rect 4934 4824 4972 4858
rect 5006 4824 5044 4858
rect 5078 4824 5116 4858
rect 5150 4824 5188 4858
rect 5222 4824 5260 4858
rect 5294 4824 5332 4858
rect 5366 4824 5404 4858
rect 5438 4824 5476 4858
rect 5510 4824 5548 4858
rect 5582 4824 5620 4858
rect 5654 4824 5692 4858
rect 5726 4824 5764 4858
rect 5798 4824 5836 4858
rect 5870 4824 5908 4858
rect 5942 4824 5980 4858
rect 6014 4824 6052 4858
rect 6086 4824 6124 4858
rect 6158 4824 6196 4858
rect 6230 4824 6268 4858
rect 6302 4824 6340 4858
rect 6374 4824 6412 4858
rect 6446 4824 6484 4858
rect 6518 4824 6556 4858
rect 6590 4824 6628 4858
rect 6662 4824 6700 4858
rect 6734 4824 6772 4858
rect 6806 4824 6844 4858
rect 6878 4824 6916 4858
rect 6950 4824 6988 4858
rect 7022 4824 7060 4858
rect 7094 4824 7132 4858
rect 7166 4824 7204 4858
rect 7238 4824 7276 4858
rect 7310 4824 7348 4858
rect 7382 4824 7420 4858
rect 7454 4824 7492 4858
rect 7526 4824 7564 4858
rect 7598 4824 7636 4858
rect 7670 4824 7708 4858
rect 7742 4824 7780 4858
rect 7814 4824 7852 4858
rect 7886 4824 7924 4858
rect 7958 4824 7996 4858
rect 8030 4824 8068 4858
rect 8102 4824 8140 4858
rect 8174 4824 8212 4858
rect 8246 4824 8284 4858
rect 8318 4824 8356 4858
rect 8390 4824 8428 4858
rect 8462 4824 8500 4858
rect 8534 4824 8572 4858
rect 8606 4824 8644 4858
rect 8678 4824 8716 4858
rect 8750 4824 8788 4858
rect 8822 4824 8860 4858
rect 8894 4824 8932 4858
rect 8966 4824 9004 4858
rect 9038 4824 9076 4858
rect 9110 4824 9148 4858
rect 9182 4824 9220 4858
rect 9254 4824 9292 4858
rect 9326 4824 9364 4858
rect 9398 4824 9436 4858
rect 9470 4824 9508 4858
rect 9542 4824 9580 4858
rect 9614 4824 9652 4858
rect 9686 4824 9724 4858
rect 9758 4824 9796 4858
rect 9830 4824 9868 4858
rect 9902 4824 9940 4858
rect 9974 4824 10012 4858
rect 10046 4824 10084 4858
rect 10118 4824 10156 4858
rect 10190 4824 10228 4858
rect 10262 4824 10300 4858
rect 10334 4824 10372 4858
rect 10406 4824 10444 4858
rect 10478 4824 10516 4858
rect 10550 4824 10588 4858
rect 10622 4824 10660 4858
rect 10694 4824 10732 4858
rect 10766 4824 10804 4858
rect 10838 4824 10876 4858
rect 10910 4824 10948 4858
rect 10982 4824 11020 4858
rect 11054 4824 11092 4858
rect 11126 4824 11164 4858
rect 11198 4824 11236 4858
rect 11270 4824 11308 4858
rect 11342 4824 11380 4858
rect 11414 4824 11452 4858
rect 11486 4824 11524 4858
rect 11558 4824 11596 4858
rect 11630 4824 11668 4858
rect 11702 4824 11740 4858
rect 11774 4824 11813 4858
rect 11847 4824 11886 4858
rect 11920 4824 11959 4858
rect 11993 4824 12032 4858
rect 12066 4824 12105 4858
rect 12139 4824 12178 4858
rect 12212 4824 12251 4858
rect 12285 4824 12324 4858
rect 12358 4824 12397 4858
rect 12431 4824 12470 4858
rect 12504 4824 12543 4858
rect 12577 4824 12616 4858
rect 12650 4824 12689 4858
rect 12723 4824 12762 4858
rect 12796 4824 12835 4858
rect 12869 4824 12908 4858
rect 12942 4824 12981 4858
rect 13015 4824 13054 4858
rect 13088 4824 13127 4858
rect 13161 4824 13200 4858
rect 13234 4824 13273 4858
rect 13307 4824 13346 4858
rect 13380 4824 13392 4858
rect -26 4818 13392 4824
rect -26 4815 35 4818
rect -26 4786 26 4815
tri 26 4787 54 4815 nw
rect -26 4779 -17 4786
rect 17 4779 26 4786
rect -26 4715 26 4727
rect -26 4651 26 4663
rect -26 4587 26 4599
tri 26 4563 51 4588 sw
rect 26 4550 13103 4563
rect 26 4543 12840 4550
rect 26 4535 333 4543
rect -26 4523 333 4535
rect 26 4471 333 4523
rect -26 4464 -17 4471
rect 17 4464 333 4471
rect -26 4459 333 4464
rect 26 4437 333 4459
rect 799 4498 12840 4543
rect 12892 4498 12906 4550
rect 12958 4498 12973 4550
rect 13025 4498 13040 4550
rect 13092 4498 13103 4550
rect 799 4486 13103 4498
rect 799 4437 12840 4486
rect 26 4434 12840 4437
rect 12892 4434 12906 4486
rect 12958 4434 12973 4486
rect 13025 4434 13040 4486
rect 13092 4434 13103 4486
rect 26 4417 13103 4434
rect -26 4395 -17 4407
rect 17 4395 26 4407
tri 26 4392 51 4417 nw
rect -26 4331 -17 4343
rect 17 4331 26 4343
rect -26 4267 -17 4279
rect 17 4267 26 4279
rect 10155 4327 10207 4333
rect 10155 4263 10207 4275
tri 10130 4233 10155 4258 se
rect -26 4210 26 4215
rect -26 4203 -17 4210
rect 17 4203 26 4210
rect 7138 4211 10155 4233
rect 7138 4205 10207 4211
rect 121 4163 265 4194
rect -26 4139 26 4151
rect 7860 4131 7906 4177
rect 9102 4131 9148 4177
rect 10098 4089 10138 4135
rect -26 4075 26 4087
rect -26 4011 26 4023
rect 7668 4013 7708 4059
rect 9237 4009 9243 4061
rect 9295 4009 9307 4061
rect 9359 4009 9365 4061
rect -26 3947 26 3959
rect 5766 3933 5806 3979
rect 5902 3933 5943 3979
tri 26 3905 51 3930 sw
rect 26 3902 10240 3905
tri 10240 3902 10243 3905 sw
tri 11368 3902 11371 3905 se
rect 11371 3902 13350 3905
rect 26 3895 10243 3902
rect -26 3888 -17 3895
rect 17 3888 10243 3895
rect -26 3883 10243 3888
rect 26 3831 10243 3883
rect -26 3819 -17 3831
rect 17 3825 10243 3831
tri 10243 3825 10320 3902 sw
tri 11291 3825 11368 3902 se
rect 11368 3901 13350 3902
rect 11368 3849 12840 3901
rect 12892 3849 12906 3901
rect 12958 3849 12973 3901
rect 13025 3849 13040 3901
rect 13092 3849 13350 3901
rect 11368 3831 13350 3849
rect 11368 3825 12840 3831
rect 17 3819 12840 3825
rect 26 3779 12840 3819
rect 12892 3779 12906 3831
rect 12958 3779 12973 3831
rect 13025 3779 13040 3831
rect 13092 3779 13350 3831
rect 26 3767 13350 3779
rect -26 3755 -17 3767
rect 17 3761 13350 3767
rect 17 3755 12840 3761
rect 26 3739 12840 3755
rect 26 3708 1516 3739
tri 1516 3708 1547 3739 nw
tri 1661 3708 1692 3739 ne
rect 1692 3709 12840 3739
rect 12892 3709 12906 3761
rect 12958 3709 12973 3761
rect 13025 3709 13040 3761
rect 13092 3709 13350 3761
rect 1692 3708 13350 3709
rect 26 3703 1511 3708
tri 1511 3703 1516 3708 nw
tri 1692 3703 1697 3708 ne
rect 1697 3703 13350 3708
rect -26 3691 -17 3703
rect 17 3691 26 3703
tri 26 3678 51 3703 nw
rect -26 3634 26 3639
rect -26 3627 -17 3634
rect 17 3627 26 3634
rect 66 3629 103 3675
rect 6875 3669 9716 3675
rect -26 3563 26 3575
rect 6927 3635 7138 3669
rect 7172 3635 7210 3669
rect 7244 3635 9454 3669
rect 9488 3635 9526 3669
rect 9560 3635 9598 3669
rect 9632 3635 9670 3669
rect 9704 3635 9716 3669
rect 6927 3629 9716 3635
rect 6875 3605 6927 3617
tri 6927 3604 6952 3629 nw
rect 7540 3595 7670 3601
rect 7540 3561 7552 3595
rect 7586 3561 7624 3595
rect 7658 3561 7670 3595
rect 7540 3555 7670 3561
rect 7882 3595 9884 3601
rect 7882 3561 7896 3595
rect 7930 3561 7968 3595
rect 8002 3561 9144 3595
rect 9178 3561 9216 3595
rect 9250 3589 9884 3595
tri 9884 3589 9896 3601 sw
rect 9250 3583 9896 3589
tri 9896 3583 9902 3589 sw
rect 9985 3583 10085 3595
rect 10137 3583 10149 3595
rect 9250 3561 9902 3583
rect 7882 3555 9902 3561
tri 9902 3555 9930 3583 sw
rect 6875 3547 6927 3553
tri 9856 3549 9862 3555 ne
rect 9862 3549 9930 3555
tri 9930 3549 9936 3555 sw
rect 9985 3549 9997 3583
rect 10031 3549 10069 3583
rect 10137 3549 10141 3583
tri 9862 3547 9864 3549 ne
rect 9864 3547 9936 3549
tri 9864 3527 9884 3547 ne
rect 9884 3527 9936 3547
tri 9936 3527 9958 3549 sw
rect 9985 3543 10085 3549
rect 10137 3543 10149 3549
rect 10201 3543 10207 3595
rect -26 3499 26 3511
rect 8247 3521 8377 3527
rect 8247 3487 8259 3521
rect 8293 3487 8331 3521
rect 8365 3487 8377 3521
rect 8247 3481 8377 3487
rect 8647 3519 9543 3527
rect 8647 3485 8659 3519
rect 8693 3485 8731 3519
rect 8765 3485 9543 3519
rect 8647 3475 9543 3485
rect 9595 3475 9607 3527
rect 9659 3475 9665 3527
tri 9884 3515 9896 3527 ne
rect 9896 3515 9958 3527
tri 9958 3515 9970 3527 sw
tri 9896 3475 9936 3515 ne
rect 9936 3475 12621 3515
tri 9936 3463 9948 3475 ne
rect 9948 3463 12621 3475
rect 12673 3463 12685 3515
rect 12737 3463 12743 3515
rect -26 3415 26 3447
rect 0 3372 10260 3379
rect 0 3194 9173 3372
rect 9279 3334 10260 3372
tri 10260 3334 10305 3379 sw
tri 10471 3334 10516 3379 se
rect 10516 3334 12778 3379
rect 9279 3194 12778 3334
rect 0 3177 12778 3194
rect -81 3109 -23 3115
rect -81 3057 -78 3109
rect -26 3057 -23 3109
tri 12750 3061 12775 3086 ne
tri 12821 3061 12846 3086 nw
tri 12906 3061 12931 3086 ne
rect -81 3045 -23 3057
rect -81 2993 -78 3045
rect -26 2993 -23 3045
rect 10897 3006 12101 3058
rect 12153 3006 12165 3058
rect 12217 3006 12223 3058
rect -81 2981 -23 2993
rect -81 2929 -78 2981
rect -26 2929 -23 2981
rect -81 2923 -23 2929
rect 0 2883 12803 2895
rect 0 2777 400 2883
rect 1010 2777 12803 2883
rect 0 2765 12803 2777
rect -81 2707 -23 2713
rect -81 2673 -69 2707
rect -35 2673 -23 2707
rect -81 2657 -23 2673
rect -81 2605 -78 2657
rect -26 2605 -23 2657
rect -81 2601 -69 2605
rect -35 2601 -23 2605
rect -81 2593 -23 2601
rect -81 2541 -78 2593
rect -26 2541 -23 2593
rect -81 2529 -69 2541
rect -35 2529 -23 2541
rect -81 2477 -78 2529
rect -26 2477 -23 2529
rect -81 2465 -69 2477
rect -35 2465 -23 2477
rect -81 2413 -78 2465
rect -26 2413 -23 2465
rect -81 2401 -69 2413
rect -35 2401 -23 2413
rect -81 2349 -78 2401
rect -26 2349 -23 2401
tri 1047 2381 1051 2385 se
rect 1051 2381 3888 2385
rect 4267 2381 4373 2385
tri 4373 2381 4377 2385 sw
tri 1041 2375 1047 2381 se
rect 1047 2375 4385 2381
rect -81 2347 -23 2349
rect -81 2313 -69 2347
rect -35 2313 -23 2347
tri 1007 2341 1041 2375 se
rect 1041 2341 1061 2375
rect 1095 2341 1134 2375
rect 1168 2341 1207 2375
rect 1241 2341 1280 2375
rect 1314 2341 1353 2375
rect 1387 2341 1426 2375
rect 1460 2341 1499 2375
rect 1533 2341 1572 2375
rect 1606 2341 1645 2375
rect 1679 2341 1718 2375
rect 1752 2341 1791 2375
rect 1825 2341 1864 2375
rect 1898 2341 1937 2375
rect 1971 2341 2010 2375
rect 2044 2341 2083 2375
rect 2117 2341 2156 2375
rect 2190 2341 2229 2375
rect 2263 2341 2302 2375
rect 2336 2341 2375 2375
rect 2409 2341 2448 2375
rect 2482 2341 2521 2375
rect 2555 2341 2594 2375
rect 2628 2341 2667 2375
rect 2701 2341 2740 2375
rect 2774 2341 2813 2375
rect 2847 2341 2886 2375
rect 2920 2341 2959 2375
rect 2993 2341 3032 2375
rect 3066 2341 3105 2375
rect 3139 2341 3178 2375
rect 3212 2341 3251 2375
rect 3285 2341 3324 2375
rect 3358 2341 3397 2375
rect 3431 2341 3470 2375
rect 3504 2341 3543 2375
rect 3577 2341 3616 2375
rect 3650 2341 3689 2375
rect 3723 2341 3762 2375
rect 3796 2341 3835 2375
rect 3869 2341 3907 2375
rect 3941 2341 3979 2375
rect 4013 2341 4051 2375
rect 4085 2341 4123 2375
rect 4157 2341 4195 2375
rect 4229 2341 4267 2375
rect 4301 2341 4339 2375
rect 4373 2341 4385 2375
tri 1001 2335 1007 2341 se
rect 1007 2335 4385 2341
tri 4385 2335 4423 2373 sw
rect -81 2307 -23 2313
tri 973 2307 1001 2335 se
rect 1001 2307 3888 2335
tri 945 2279 973 2307 se
rect 973 2279 3888 2307
rect 700 2255 3888 2279
rect 4267 2279 4423 2335
tri 4423 2279 4479 2335 sw
rect 9524 2307 9543 2359
rect 9595 2307 9607 2359
rect 9659 2307 9665 2359
rect 9781 2307 9827 2353
tri 12988 2282 13013 2307 ne
rect 4267 2255 12909 2279
rect 700 2149 3023 2255
tri 3027 2149 3133 2255 nw
tri 4267 2149 4373 2255 ne
rect 4373 2149 12909 2255
rect -75 2014 26 2042
rect -75 1962 -26 2014
rect -75 1950 26 1962
rect -75 1898 -26 1950
rect -75 1886 26 1898
rect -75 1834 -26 1886
rect -75 1822 26 1834
rect -75 1770 -26 1822
rect -75 1758 26 1770
rect -75 1706 -26 1758
tri 742 1753 743 1754 se
rect 743 1753 13369 1754
tri 731 1742 742 1753 se
rect 742 1752 13369 1753
rect 742 1742 12837 1752
tri 718 1729 731 1742 se
rect 731 1729 12557 1742
tri 712 1723 718 1729 se
rect 718 1723 12557 1729
rect -75 1694 26 1706
rect -75 1642 -26 1694
tri 678 1689 712 1723 se
rect 712 1689 9155 1723
rect 9189 1689 9227 1723
rect 9261 1708 12557 1723
rect 12591 1708 12837 1742
rect 9261 1700 12837 1708
rect 12889 1700 12904 1752
rect 12956 1700 12971 1752
rect 13023 1700 13038 1752
rect 13090 1700 13105 1752
rect 13157 1700 13172 1752
rect 13224 1700 13239 1752
rect 13291 1700 13306 1752
rect 13358 1700 13369 1752
rect 9261 1689 13369 1700
tri 672 1683 678 1689 se
rect 678 1683 13369 1689
tri 659 1670 672 1683 se
rect 672 1680 13369 1683
rect 672 1670 12837 1680
tri 642 1653 659 1670 se
rect 659 1653 12557 1670
rect -75 1636 26 1642
tri 26 1636 43 1653 sw
tri 625 1636 642 1653 se
rect 642 1636 12557 1653
rect 12591 1636 12837 1670
rect -75 1630 43 1636
rect -75 1578 -26 1630
rect 26 1598 43 1630
tri 43 1598 81 1636 sw
tri 587 1598 625 1636 se
rect 625 1628 12837 1636
rect 12889 1628 12904 1680
rect 12956 1628 12971 1680
rect 13023 1628 13038 1680
rect 13090 1628 13105 1680
rect 13157 1628 13172 1680
rect 13224 1628 13239 1680
rect 13291 1628 13306 1680
rect 13358 1628 13369 1680
rect 625 1608 13369 1628
rect 625 1598 12837 1608
rect 26 1578 81 1598
rect -75 1566 81 1578
rect -75 1514 -26 1566
rect 26 1564 81 1566
tri 81 1564 115 1598 sw
tri 553 1564 587 1598 se
rect 587 1564 12557 1598
rect 12591 1564 12837 1598
rect 26 1514 115 1564
rect -75 1502 115 1514
rect -75 1450 -26 1502
rect 26 1488 115 1502
tri 115 1488 191 1564 sw
tri 544 1555 553 1564 se
rect 553 1556 12837 1564
rect 12889 1556 12904 1608
rect 12956 1556 12971 1608
rect 13023 1556 13038 1608
rect 13090 1556 13105 1608
rect 13157 1556 13172 1608
rect 13224 1556 13239 1608
rect 13291 1556 13306 1608
rect 13358 1556 13369 1608
rect 553 1555 13369 1556
tri 477 1488 544 1555 se
rect 544 1552 13369 1555
rect 544 1488 900 1552
tri 900 1488 964 1552 nw
rect 26 1474 886 1488
tri 886 1474 900 1488 nw
rect 26 1450 852 1474
rect -75 1440 852 1450
tri 852 1440 886 1474 nw
rect -75 1438 814 1440
rect -75 1386 -26 1438
rect 26 1402 814 1438
tri 814 1402 852 1440 nw
rect 9468 1403 9505 1480
rect 12551 1474 12597 1486
rect 12551 1440 12557 1474
rect 12591 1440 12597 1474
rect 12551 1402 12597 1440
rect 26 1386 781 1402
rect -75 1374 781 1386
rect -75 1322 -26 1374
rect 26 1322 781 1374
tri 781 1369 814 1402 nw
rect -75 1179 781 1322
rect 12551 1368 12557 1402
rect 12591 1368 12597 1402
rect 12551 1330 12597 1368
rect 12551 1296 12557 1330
rect 12591 1296 12597 1330
rect 12551 1284 12597 1296
rect -75 1145 66 1179
rect 100 1145 141 1179
rect 175 1145 216 1179
rect 250 1145 291 1179
rect 325 1145 367 1179
rect 401 1145 443 1179
rect 477 1145 519 1179
rect 553 1145 595 1179
rect 629 1145 781 1179
rect -75 1107 781 1145
rect -75 1073 66 1107
rect 100 1073 141 1107
rect 175 1073 216 1107
rect 250 1073 291 1107
rect 325 1073 367 1107
rect 401 1073 443 1107
rect 477 1073 519 1107
rect 553 1073 595 1107
rect 629 1073 781 1107
rect -75 1035 781 1073
rect -75 1001 66 1035
rect 100 1001 141 1035
rect 175 1001 216 1035
rect 250 1001 291 1035
rect 325 1001 367 1035
rect 401 1001 443 1035
rect 477 1001 519 1035
rect 553 1001 595 1035
rect 629 1001 781 1035
rect 857 1221 12908 1228
rect 857 1043 8463 1221
rect 8713 1043 12908 1221
rect 857 1026 12908 1043
rect -75 963 781 1001
rect -75 929 66 963
rect 100 929 141 963
rect 175 929 216 963
rect 250 929 291 963
rect 325 929 367 963
rect 401 929 443 963
rect 477 929 519 963
rect 553 929 595 963
rect 629 929 781 963
rect -75 910 781 929
tri 781 910 824 953 sw
rect -75 898 824 910
tri 824 898 836 910 sw
tri 12546 898 12558 910 se
rect 12558 898 12604 910
rect -75 891 836 898
rect -75 857 66 891
rect 100 857 141 891
rect 175 857 216 891
rect 250 857 291 891
rect 325 857 367 891
rect 401 857 443 891
rect 477 857 519 891
rect 553 857 595 891
rect 629 864 836 891
tri 836 864 870 898 sw
tri 12512 864 12546 898 se
rect 12546 864 12564 898
rect 12598 864 12604 898
rect 629 858 870 864
tri 870 858 876 864 sw
tri 12506 858 12512 864 se
rect 12512 858 12604 864
rect 629 857 876 858
rect -75 851 876 857
tri 876 851 883 858 sw
tri 12138 851 12145 858 se
rect 12145 851 12604 858
rect -75 839 883 851
tri 883 839 895 851 sw
tri 12126 839 12138 851 se
rect 12138 839 12604 851
tri -75 826 -62 839 ne
rect -62 826 895 839
tri 895 826 908 839 sw
tri 12113 826 12126 839 se
rect 12126 826 12604 839
tri -62 813 -49 826 ne
rect -49 813 12564 826
tri -49 781 -17 813 ne
rect -17 781 12190 813
tri -17 747 17 781 ne
rect 17 747 121 781
rect 155 747 193 781
rect 227 747 265 781
rect 299 747 337 781
rect 371 747 409 781
rect 443 747 481 781
rect 515 747 553 781
rect 587 747 625 781
rect 659 747 697 781
rect 731 747 769 781
rect 803 747 841 781
rect 875 747 913 781
rect 947 747 985 781
rect 1019 747 1057 781
rect 1091 747 1129 781
rect 1163 747 1201 781
rect 1235 747 1273 781
rect 1307 747 1345 781
rect 1379 747 1417 781
rect 1451 747 1489 781
rect 1523 747 1561 781
rect 1595 747 1633 781
rect 1667 747 1705 781
rect 1739 747 1777 781
rect 1811 747 1849 781
rect 1883 747 1921 781
rect 1955 747 1993 781
rect 2027 747 2065 781
rect 2099 747 2137 781
rect 2171 747 2209 781
rect 2243 747 2281 781
rect 2315 747 2353 781
rect 2387 747 2425 781
rect 2459 747 2497 781
rect 2531 747 2569 781
rect 2603 747 2641 781
rect 2675 747 2713 781
rect 2747 747 2785 781
rect 2819 747 2857 781
rect 2891 747 2929 781
rect 2963 747 3001 781
rect 3035 747 3073 781
rect 3107 747 3145 781
rect 3179 747 3217 781
rect 3251 747 3289 781
rect 3323 747 3361 781
rect 3395 747 3433 781
rect 3467 747 3505 781
rect 3539 747 3577 781
rect 3611 747 3649 781
rect 3683 747 3721 781
rect 3755 747 3793 781
rect 3827 747 3865 781
rect 3899 747 3937 781
rect 3971 747 4009 781
rect 4043 747 4081 781
rect 4115 747 4153 781
rect 4187 747 4225 781
rect 4259 747 4297 781
rect 4331 747 4369 781
rect 4403 747 4441 781
rect 4475 747 4513 781
rect 4547 747 4585 781
rect 4619 747 4657 781
rect 4691 747 4729 781
rect 4763 747 4801 781
rect 4835 747 4873 781
rect 4907 747 4945 781
rect 4979 747 5017 781
rect 5051 747 5089 781
rect 5123 747 5161 781
rect 5195 747 5233 781
rect 5267 747 5305 781
rect 5339 747 5377 781
rect 5411 747 5449 781
rect 5483 747 5521 781
rect 5555 747 5593 781
rect 5627 747 5665 781
rect 5699 747 5737 781
rect 5771 747 5809 781
rect 5843 747 5881 781
rect 5915 747 5953 781
rect 5987 747 6025 781
rect 6059 747 6097 781
rect 6131 747 6169 781
rect 6203 747 6241 781
rect 6275 747 6313 781
rect 6347 747 6385 781
rect 6419 747 6457 781
rect 6491 747 6529 781
rect 6563 747 6601 781
rect 6635 747 6673 781
rect 6707 747 6745 781
rect 6779 747 6817 781
rect 6851 747 6889 781
rect 6923 747 6961 781
rect 6995 747 7033 781
rect 7067 747 7105 781
rect 7139 747 7177 781
rect 7211 747 7249 781
rect 7283 747 7321 781
rect 7355 747 7393 781
rect 7427 747 7465 781
rect 7499 747 7537 781
rect 7571 747 7609 781
rect 7643 747 7681 781
rect 7715 747 7753 781
rect 7787 747 7825 781
rect 7859 747 7897 781
rect 7931 747 7969 781
rect 8003 747 8041 781
rect 8075 747 8113 781
rect 8147 747 8185 781
rect 8219 747 8257 781
rect 8291 747 8329 781
rect 8363 747 8401 781
rect 8435 747 8473 781
rect 8507 747 8545 781
rect 8579 747 8617 781
rect 8651 747 8689 781
rect 8723 747 8761 781
rect 8795 747 8833 781
rect 8867 747 8905 781
rect 8939 747 8977 781
rect 9011 747 9049 781
rect 9083 747 9121 781
rect 9155 747 9193 781
rect 9227 747 9265 781
rect 9299 747 9337 781
rect 9371 747 9409 781
rect 9443 747 9481 781
rect 9515 747 9553 781
rect 9587 747 9625 781
rect 9659 747 9697 781
rect 9731 747 9769 781
rect 9803 747 9841 781
rect 9875 747 9913 781
rect 9947 747 9985 781
rect 10019 747 10057 781
rect 10091 747 10129 781
rect 10163 747 10201 781
rect 10235 747 10273 781
rect 10307 747 10345 781
rect 10379 747 10417 781
rect 10451 747 10489 781
rect 10523 747 10561 781
rect 10595 747 10633 781
rect 10667 747 10705 781
rect 10739 747 10777 781
rect 10811 747 10849 781
rect 10883 747 10921 781
rect 10955 747 10993 781
rect 11027 747 11065 781
rect 11099 747 11137 781
rect 11171 747 11209 781
rect 11243 747 11281 781
rect 11315 747 11353 781
rect 11387 747 11425 781
rect 11459 747 11497 781
rect 11531 747 11569 781
rect 11603 747 11641 781
rect 11675 747 11713 781
rect 11747 747 11785 781
rect 11819 747 11857 781
rect 11891 747 11929 781
rect 11963 747 12001 781
rect 12035 747 12073 781
rect 12107 779 12190 781
rect 12224 779 12262 813
rect 12296 779 12334 813
rect 12368 779 12406 813
rect 12440 779 12478 813
rect 12512 792 12564 813
rect 12598 792 12604 826
rect 12512 779 12604 792
rect 12107 747 12604 779
tri 17 743 21 747 ne
rect 21 734 12604 747
rect 21 702 12269 734
tri 12269 702 12301 734 nw
<< via1 >>
rect -26 4752 -17 4779
rect -17 4752 17 4779
rect 17 4752 26 4779
rect -26 4727 26 4752
rect -26 4714 26 4715
rect -26 4680 -17 4714
rect -17 4680 17 4714
rect 17 4680 26 4714
rect -26 4663 26 4680
rect -26 4642 26 4651
rect -26 4608 -17 4642
rect -17 4608 17 4642
rect 17 4608 26 4642
rect -26 4599 26 4608
rect -26 4570 26 4587
rect -26 4536 -17 4570
rect -17 4536 17 4570
rect 17 4536 26 4570
rect -26 4535 26 4536
rect -26 4498 26 4523
rect -26 4471 -17 4498
rect -17 4471 17 4498
rect 17 4471 26 4498
rect -26 4426 26 4459
rect 12840 4498 12892 4550
rect 12906 4498 12958 4550
rect 12973 4498 13025 4550
rect 13040 4498 13092 4550
rect 12840 4434 12892 4486
rect 12906 4434 12958 4486
rect 12973 4434 13025 4486
rect 13040 4434 13092 4486
rect -26 4407 -17 4426
rect -17 4407 17 4426
rect 17 4407 26 4426
rect -26 4392 -17 4395
rect -17 4392 17 4395
rect 17 4392 26 4395
rect -26 4354 26 4392
rect -26 4343 -17 4354
rect -17 4343 17 4354
rect 17 4343 26 4354
rect -26 4320 -17 4331
rect -17 4320 17 4331
rect 17 4320 26 4331
rect -26 4282 26 4320
rect -26 4279 -17 4282
rect -17 4279 17 4282
rect 17 4279 26 4282
rect -26 4248 -17 4267
rect -17 4248 17 4267
rect 17 4248 26 4267
rect 10155 4275 10207 4327
rect -26 4215 26 4248
rect 10155 4211 10207 4263
rect -26 4176 -17 4203
rect -17 4176 17 4203
rect 17 4176 26 4203
rect -26 4151 26 4176
rect -26 4138 26 4139
rect -26 4104 -17 4138
rect -17 4104 17 4138
rect 17 4104 26 4138
rect -26 4087 26 4104
rect -26 4066 26 4075
rect -26 4032 -17 4066
rect -17 4032 17 4066
rect 17 4032 26 4066
rect -26 4023 26 4032
rect -26 3994 26 4011
rect 9243 4009 9295 4061
rect 9307 4009 9359 4061
rect -26 3960 -17 3994
rect -17 3960 17 3994
rect 17 3960 26 3994
rect -26 3959 26 3960
rect -26 3922 26 3947
rect -26 3895 -17 3922
rect -17 3895 17 3922
rect 17 3895 26 3922
rect -26 3850 26 3883
rect -26 3831 -17 3850
rect -17 3831 17 3850
rect 17 3831 26 3850
rect 12840 3849 12892 3901
rect 12906 3849 12958 3901
rect 12973 3849 13025 3901
rect 13040 3849 13092 3901
rect -26 3816 -17 3819
rect -17 3816 17 3819
rect 17 3816 26 3819
rect -26 3778 26 3816
rect 12840 3779 12892 3831
rect 12906 3779 12958 3831
rect 12973 3779 13025 3831
rect 13040 3779 13092 3831
rect -26 3767 -17 3778
rect -17 3767 17 3778
rect 17 3767 26 3778
rect -26 3744 -17 3755
rect -17 3744 17 3755
rect 17 3744 26 3755
rect -26 3706 26 3744
rect 12840 3709 12892 3761
rect 12906 3709 12958 3761
rect 12973 3709 13025 3761
rect 13040 3709 13092 3761
rect -26 3703 -17 3706
rect -17 3703 17 3706
rect 17 3703 26 3706
rect -26 3672 -17 3691
rect -17 3672 17 3691
rect 17 3672 26 3691
rect -26 3639 26 3672
rect -26 3600 -17 3627
rect -17 3600 17 3627
rect 17 3600 26 3627
rect -26 3575 26 3600
rect -26 3562 26 3563
rect -26 3528 -17 3562
rect -17 3528 17 3562
rect 17 3528 26 3562
rect 6875 3617 6927 3669
rect 6875 3553 6927 3605
rect 10085 3583 10137 3595
rect 10149 3583 10201 3595
rect 10085 3549 10103 3583
rect 10103 3549 10137 3583
rect 10149 3549 10175 3583
rect 10175 3549 10201 3583
rect -26 3511 26 3528
rect 10085 3543 10137 3549
rect 10149 3543 10201 3549
rect -26 3490 26 3499
rect -26 3456 -17 3490
rect -17 3456 17 3490
rect 17 3456 26 3490
rect 9543 3475 9595 3527
rect 9607 3475 9659 3527
rect 12621 3463 12673 3515
rect 12685 3463 12737 3515
rect -26 3447 26 3456
rect -78 3108 -26 3109
rect -78 3074 -69 3108
rect -69 3074 -35 3108
rect -35 3074 -26 3108
rect -78 3057 -26 3074
rect -78 3036 -26 3045
rect -78 3002 -69 3036
rect -69 3002 -35 3036
rect -35 3002 -26 3036
rect -78 2993 -26 3002
rect 12101 3006 12153 3058
rect 12165 3006 12217 3058
rect -78 2964 -26 2981
rect -78 2930 -69 2964
rect -69 2930 -35 2964
rect -35 2930 -26 2964
rect -78 2929 -26 2930
rect -78 2635 -26 2657
rect -78 2605 -69 2635
rect -69 2605 -35 2635
rect -35 2605 -26 2635
rect -78 2563 -26 2593
rect -78 2541 -69 2563
rect -69 2541 -35 2563
rect -35 2541 -26 2563
rect -78 2491 -26 2529
rect -78 2477 -69 2491
rect -69 2477 -35 2491
rect -35 2477 -26 2491
rect -78 2457 -69 2465
rect -69 2457 -35 2465
rect -35 2457 -26 2465
rect -78 2419 -26 2457
rect -78 2413 -69 2419
rect -69 2413 -35 2419
rect -35 2413 -26 2419
rect -78 2385 -69 2401
rect -69 2385 -35 2401
rect -35 2385 -26 2401
rect -78 2349 -26 2385
rect 9543 2307 9595 2359
rect 9607 2307 9659 2359
rect -26 1962 26 2014
rect -26 1898 26 1950
rect -26 1834 26 1886
rect -26 1770 26 1822
rect -26 1706 26 1758
rect -26 1642 26 1694
rect 12837 1700 12889 1752
rect 12904 1700 12956 1752
rect 12971 1700 13023 1752
rect 13038 1700 13090 1752
rect 13105 1700 13157 1752
rect 13172 1700 13224 1752
rect 13239 1700 13291 1752
rect 13306 1700 13358 1752
rect -26 1578 26 1630
rect 12837 1628 12889 1680
rect 12904 1628 12956 1680
rect 12971 1628 13023 1680
rect 13038 1628 13090 1680
rect 13105 1628 13157 1680
rect 13172 1628 13224 1680
rect 13239 1628 13291 1680
rect 13306 1628 13358 1680
rect -26 1514 26 1566
rect -26 1450 26 1502
rect 12837 1556 12889 1608
rect 12904 1556 12956 1608
rect 12971 1556 13023 1608
rect 13038 1556 13090 1608
rect 13105 1556 13157 1608
rect 13172 1556 13224 1608
rect 13239 1556 13291 1608
rect 13306 1556 13358 1608
rect -26 1386 26 1438
rect -26 1322 26 1374
<< metal2 >>
rect -26 4779 26 4785
rect -26 4715 26 4727
rect -26 4651 26 4663
rect -26 4587 26 4599
rect -26 4523 26 4535
rect -26 4459 26 4471
rect -26 4395 26 4407
rect -26 4331 26 4343
rect 12828 4550 13101 4564
rect 12828 4498 12840 4550
rect 12892 4498 12906 4550
rect 12958 4498 12973 4550
rect 13025 4498 13040 4550
rect 13092 4498 13101 4550
rect 12828 4486 13101 4498
rect 12828 4434 12840 4486
rect 12892 4434 12906 4486
rect 12958 4434 12973 4486
rect 13025 4434 13040 4486
rect 13092 4434 13101 4486
rect -26 4267 26 4279
rect -26 4203 26 4215
rect -26 4139 26 4151
rect -26 4075 26 4087
rect 10155 4327 10207 4333
rect 10155 4263 10207 4275
rect -26 4011 26 4023
rect 9237 4009 9243 4061
rect 9295 4009 9307 4061
rect 9359 4009 9365 4061
rect -26 3947 26 3959
rect -26 3883 26 3895
rect -26 3819 26 3831
rect -26 3755 26 3767
rect -26 3691 26 3703
rect -26 3627 26 3639
rect -26 3563 26 3575
rect 6875 3669 6927 3675
rect 6875 3605 6927 3617
rect 6875 3535 6927 3553
rect 9313 3527 9365 4009
tri 10130 3595 10155 3620 se
rect 10155 3595 10207 4211
rect 12828 3901 13101 4434
rect 12828 3849 12840 3901
rect 12892 3849 12906 3901
rect 12958 3849 12973 3901
rect 13025 3849 13040 3901
rect 13092 3849 13101 3901
rect 12828 3831 13101 3849
rect 12828 3779 12840 3831
rect 12892 3779 12906 3831
rect 12958 3779 12973 3831
rect 13025 3779 13040 3831
rect 13092 3779 13101 3831
rect 12828 3761 13101 3779
rect 12828 3709 12840 3761
rect 12892 3709 12906 3761
rect 12958 3709 12973 3761
rect 13025 3709 13040 3761
rect 13092 3709 13101 3761
rect 10324 3623 10382 3675
rect 10079 3543 10085 3595
rect 10137 3543 10149 3595
rect 10201 3543 10207 3595
rect -26 3499 26 3511
tri -78 3115 -26 3167 se
rect -26 3115 26 3447
rect -78 3109 26 3115
rect -26 3057 26 3109
rect -78 3045 26 3057
rect -26 2993 26 3045
rect -78 2981 26 2993
rect -26 2929 26 2981
rect -78 2923 26 2929
tri -78 2871 -26 2923 ne
tri -78 2663 -26 2715 se
rect -26 2663 26 2923
rect 9537 3475 9543 3527
rect 9595 3475 9607 3527
rect 9659 3475 9665 3527
rect -78 2657 26 2663
rect -26 2605 26 2657
rect -78 2593 26 2605
rect -26 2541 26 2593
rect 7368 2564 7411 2715
rect -78 2529 26 2541
rect -26 2477 26 2529
rect -78 2465 26 2477
rect -26 2413 26 2465
rect -78 2401 26 2413
rect -26 2349 26 2401
rect -78 2343 26 2349
tri -78 2307 -42 2343 ne
rect -42 2307 26 2343
rect 9537 2359 9665 3475
rect 12615 3463 12621 3515
rect 12673 3463 12685 3515
rect 12737 3463 12743 3515
rect 12095 3006 12101 3058
rect 12153 3006 12165 3058
rect 12217 3006 12223 3058
rect 9537 2307 9543 2359
rect 9595 2307 9607 2359
rect 9659 2307 9665 2359
tri -42 2291 -26 2307 ne
rect -26 2014 26 2307
rect -26 1950 26 1962
rect 9855 1940 9902 1992
rect -26 1886 26 1898
rect -26 1822 26 1834
rect 12828 1789 13101 3709
rect -26 1758 26 1770
rect -26 1694 26 1706
rect -26 1630 26 1642
rect -26 1566 26 1578
rect 12831 1752 13364 1753
rect 12831 1700 12837 1752
rect 12889 1700 12904 1752
rect 12956 1700 12971 1752
rect 13023 1700 13038 1752
rect 13090 1700 13105 1752
rect 13157 1700 13172 1752
rect 13224 1700 13239 1752
rect 13291 1700 13306 1752
rect 13358 1700 13364 1752
rect 12831 1680 13364 1700
rect 12831 1628 12837 1680
rect 12889 1628 12904 1680
rect 12956 1628 12971 1680
rect 13023 1628 13038 1680
rect 13090 1628 13105 1680
rect 13157 1628 13172 1680
rect 13224 1628 13239 1680
rect 13291 1628 13306 1680
rect 13358 1628 13364 1680
rect 12831 1608 13364 1628
rect 12831 1556 12837 1608
rect 12889 1556 12904 1608
rect 12956 1556 12971 1608
rect 13023 1556 13038 1608
rect 13090 1556 13105 1608
rect 13157 1556 13172 1608
rect 13224 1556 13239 1608
rect 13291 1556 13306 1608
rect 13358 1556 13364 1608
rect 12831 1555 13364 1556
rect -26 1502 26 1514
rect -26 1438 26 1450
rect -26 1374 26 1386
rect -26 1316 26 1322
use sky130_fd_pr__via_l1m1__example_55959141808269  sky130_fd_pr__via_l1m1__example_55959141808269_0
timestamp 1633016201
transform 0 -1 17 1 0 3456
box 0 0 1 1
use sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos  sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos_0
timestamp 1633016201
transform 1 0 660 0 1 906
box -162 -119 12773 3859
use sky130_fd_pr__via_l1m1__example_55959141808266  sky130_fd_pr__via_l1m1__example_55959141808266_0
timestamp 1633016201
transform -1 0 8713 0 -1 1221
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808267  sky130_fd_pr__via_l1m1__example_55959141808267_0
timestamp 1633016201
transform 0 -1 799 -1 0 4543
box 0 0 1 1
use sky130_fd_io__feas_com_pupredrvr_weak  sky130_fd_io__feas_com_pupredrvr_weak_0
timestamp 1633016201
transform -1 0 7791 0 1 2798
box 21 7 731 1967
use sky130_fd_io__com_pdpredrvr_weak  sky130_fd_io__com_pdpredrvr_weak_0
timestamp 1633016201
transform -1 0 8515 0 1 2797
box -85 8 809 1568
use sky130_fd_io__com_pupredrvr_strong_slow  sky130_fd_io__com_pupredrvr_strong_slow_0
timestamp 1633016201
transform -1 0 10215 0 1 2797
box -85 0 913 1568
use sky130_fd_io__com_pdpredrvr_strong_slow  sky130_fd_io__com_pdpredrvr_strong_slow_0
timestamp 1633016201
transform -1 0 9387 0 1 2797
box 0 0 872 1568
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_0
timestamp 1633016201
transform 1 0 9173 0 -1 3372
box 0 0 1 1
use sky130_fd_io__gpio_ovtv2_pupredrvr_strong  sky130_fd_io__gpio_ovtv2_pupredrvr_strong_0
timestamp 1633016201
transform 1 0 66 0 1 2133
box -66 -59 7278 2632
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1633016201
transform 1 0 -69 0 -1 3108
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808270  sky130_fd_pr__via_l1m1__example_55959141808270_0
timestamp 1633016201
transform 1 0 55 0 1 4824
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_0
timestamp 1633016201
transform 1 0 9454 0 1 3635
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1633016201
transform 0 1 12557 -1 0 1474
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1633016201
transform 0 -1 12591 1 0 1564
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1633016201
transform -1 0 10175 0 1 3549
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808261  sky130_fd_pr__via_m1m2__example_55959141808261_0
timestamp 1633016201
transform 0 -1 -26 1 0 2923
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1633016201
transform 1 0 9537 0 1 2307
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1633016201
transform -1 0 9665 0 -1 3527
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1633016201
transform 1 0 12615 0 1 3463
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1633016201
transform -1 0 9365 0 -1 4061
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1633016201
transform 1 0 10079 0 -1 3595
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1633016201
transform 0 -1 10207 -1 0 4333
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1633016201
transform 0 1 6875 1 0 3547
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1633016201
transform 1 0 8659 0 1 3485
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1633016201
transform -1 0 8002 0 1 3561
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1633016201
transform -1 0 9250 0 1 3561
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1633016201
transform 1 0 7138 0 1 3635
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808268  sky130_fd_pr__via_l1m1__example_55959141808268_0
timestamp 1633016201
transform 1 0 -69 0 -1 2707
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808265  sky130_fd_pr__via_l1m1__example_55959141808265_0
timestamp 1633016201
transform 0 1 400 -1 0 2883
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808263  sky130_fd_pr__via_m1m2__example_55959141808263_0
timestamp 1633016201
transform 0 -1 26 -1 0 2020
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808262  sky130_fd_pr__via_m1m2__example_55959141808262_0
timestamp 1633016201
transform 0 -1 26 -1 0 4785
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808259  sky130_fd_pr__via_m1m2__example_55959141808259_0
timestamp 1633016201
transform 0 -1 -26 -1 0 2663
box 0 0 1 1
<< labels >>
flabel metal2 s 10324 3623 10382 3675 3 FreeSans 300 0 0 0 PD_H[3]
port 1 nsew
flabel metal2 s 9855 1940 9902 1992 3 FreeSans 300 180 0 0 PD_H[2]
port 2 nsew
flabel metal2 s 7368 2564 7411 2715 3 FreeSans 520 0 0 0 PDEN_H_N[1]
port 3 nsew
flabel metal2 s 6875 3535 6927 3587 3 FreeSans 300 0 0 0 DRVHI_H
port 4 nsew
flabel metal2 s 12696 3463 12743 3515 7 FreeSans 300 180 0 0 DRVLO_H_N
port 5 nsew
flabel metal1 s 9468 1403 9505 1480 3 FreeSans 520 90 0 0 NSW_EN
port 6 nsew
flabel metal1 s 9539 2307 9587 2353 3 FreeSans 520 90 0 0 EN_CMOS_B
port 7 nsew
flabel metal1 s 5902 3933 5943 3979 3 FreeSans 300 0 0 0 PU_H_N[3]
port 8 nsew
flabel metal1 s 5766 3933 5806 3979 7 FreeSans 300 0 0 0 PU_H_N[2]
port 9 nsew
flabel metal1 s 10098 4089 10138 4135 3 FreeSans 300 0 0 0 PU_H_N[1]
port 10 nsew
flabel metal1 s 7668 4013 7708 4059 3 FreeSans 300 0 0 0 PU_H_N[0]
port 11 nsew
flabel metal1 s 9102 4131 9148 4177 3 FreeSans 300 0 0 0 PD_H[1]
port 12 nsew
flabel metal1 s 7860 4131 7906 4177 3 FreeSans 300 0 0 0 PD_H[0]
port 13 nsew
flabel metal1 s 9781 2307 9827 2353 3 FreeSans 300 0 0 0 SLOW_H
port 14 nsew
flabel metal1 s 121 4163 265 4194 3 FreeSans 520 0 0 0 PUEN_H[1]
port 15 nsew
flabel metal1 s 7550 3563 7644 3594 3 FreeSans 520 0 0 0 PUEN_H[0]
port 16 nsew
flabel metal1 s 8276 3492 8362 3516 3 FreeSans 520 0 0 0 PDEN_H_N[0]
port 17 nsew
flabel metal1 s 12736 3177 12778 3379 7 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 12866 3703 12908 3905 7 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 12871 4417 12908 4563 7 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 12760 2765 12802 2895 7 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 12866 2149 12908 2279 7 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 12866 1026 12908 1228 7 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 12866 1552 12908 1754 7 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 43 1128 85 1258 3 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 935 1026 977 1228 3 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 1112 2149 1154 2279 3 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 0 2765 42 2895 3 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 0 4417 37 4563 3 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 0 3703 42 3905 3 FreeSans 300 0 0 0 VCC_IO
port 19 nsew
flabel metal1 s 0 3177 42 3379 3 FreeSans 300 0 0 0 VGND_IO
port 18 nsew
flabel metal1 s 66 3629 103 3675 7 FreeSans 300 180 0 0 SLOW_H_N
port 20 nsew
flabel comment s 10763 779 10763 779 0 FreeSans 440 0 0 0 LIJUMPER_OK
flabel comment s 4 2252 4 2252 0 FreeSans 440 270 0 0 LIJUMPER_OK
flabel comment s 353 2539 353 2539 0 FreeSans 300 90 0 0 CONDIODE
flabel comment s 10244 3956 10244 3956 0 FreeSans 300 0 0 0 PDEN_H_N1
flabel comment s 9376 4044 9376 4044 0 FreeSans 300 0 0 0 PDEN_H_N1
flabel comment s 7497 3968 7497 3968 0 FreeSans 300 0 0 0 PDEN_H_N1
flabel comment s 7988 3576 7988 3576 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 9129 3579 9129 3579 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 10392 3490 10392 3490 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 8484 4228 8484 4228 0 FreeSans 300 0 0 0 PUEN_H1
flabel comment s 9328 4228 9328 4228 0 FreeSans 300 0 0 0 PUEN_H1
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 37174608
string GDS_START 37082662
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1310 -3013 14114 1268
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_1
timestamp 1633016201
transform 1 0 12853 0 1 -1753
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_0
timestamp 1633016201
transform 1 0 -50 0 1 7
box 0 0 1 1
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 27771720
string GDS_START 27768568
<< end >>

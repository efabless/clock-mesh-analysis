magic
tech sky130A
magscale 1 2
timestamp 1633016303
<< checkpaint >>
rect -1326 -1303 1806 2157
<< nwell >>
rect -66 377 546 897
<< pwell >>
rect 54 43 476 292
rect -26 -43 506 43
<< mvnmos >>
rect 137 116 237 266
rect 293 116 393 266
<< mvpmos >>
rect 137 443 237 743
rect 293 443 393 743
<< mvndiff >>
rect 80 258 137 266
rect 80 224 92 258
rect 126 224 137 258
rect 80 158 137 224
rect 80 124 92 158
rect 126 124 137 158
rect 80 116 137 124
rect 237 258 293 266
rect 237 224 248 258
rect 282 224 293 258
rect 237 158 293 224
rect 237 124 248 158
rect 282 124 293 158
rect 237 116 293 124
rect 393 258 450 266
rect 393 224 404 258
rect 438 224 450 258
rect 393 158 450 224
rect 393 124 404 158
rect 438 124 450 158
rect 393 116 450 124
<< mvpdiff >>
rect 80 735 137 743
rect 80 701 92 735
rect 126 701 137 735
rect 80 652 137 701
rect 80 618 92 652
rect 126 618 137 652
rect 80 568 137 618
rect 80 534 92 568
rect 126 534 137 568
rect 80 485 137 534
rect 80 451 92 485
rect 126 451 137 485
rect 80 443 137 451
rect 237 735 293 743
rect 237 701 248 735
rect 282 701 293 735
rect 237 652 293 701
rect 237 618 248 652
rect 282 618 293 652
rect 237 568 293 618
rect 237 534 248 568
rect 282 534 293 568
rect 237 485 293 534
rect 237 451 248 485
rect 282 451 293 485
rect 237 443 293 451
rect 393 735 450 743
rect 393 701 404 735
rect 438 701 450 735
rect 393 652 450 701
rect 393 618 404 652
rect 438 618 450 652
rect 393 568 450 618
rect 393 534 404 568
rect 438 534 450 568
rect 393 485 450 534
rect 393 451 404 485
rect 438 451 450 485
rect 393 443 450 451
<< mvndiffc >>
rect 92 224 126 258
rect 92 124 126 158
rect 248 224 282 258
rect 248 124 282 158
rect 404 224 438 258
rect 404 124 438 158
<< mvpdiffc >>
rect 92 701 126 735
rect 92 618 126 652
rect 92 534 126 568
rect 92 451 126 485
rect 248 701 282 735
rect 248 618 282 652
rect 248 534 282 568
rect 248 451 282 485
rect 404 701 438 735
rect 404 618 438 652
rect 404 534 438 568
rect 404 451 438 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
<< poly >>
rect 137 743 237 769
rect 293 743 393 769
rect 137 417 237 443
rect 293 417 393 443
rect 137 376 393 417
rect 80 360 393 376
rect 80 326 96 360
rect 130 326 164 360
rect 198 326 393 360
rect 80 310 393 326
rect 137 292 393 310
rect 137 266 237 292
rect 293 266 393 292
rect 137 90 237 116
rect 293 90 393 116
<< polycont >>
rect 96 326 130 360
rect 164 326 198 360
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 22 735 212 751
rect 22 701 28 735
rect 62 701 92 735
rect 134 701 172 735
rect 206 701 212 735
rect 22 652 212 701
rect 22 618 92 652
rect 126 618 212 652
rect 22 568 212 618
rect 22 534 92 568
rect 126 534 212 568
rect 22 485 212 534
rect 22 451 92 485
rect 126 451 212 485
rect 22 435 212 451
rect 248 735 298 751
rect 282 701 298 735
rect 248 652 298 701
rect 282 618 298 652
rect 248 568 298 618
rect 282 534 298 568
rect 248 485 298 534
rect 282 451 298 485
rect 25 360 214 376
rect 25 326 96 360
rect 130 326 164 360
rect 198 326 214 360
rect 25 310 214 326
rect 248 356 298 451
rect 336 735 454 751
rect 336 701 342 735
rect 376 701 404 735
rect 448 701 454 735
rect 336 652 454 701
rect 336 618 404 652
rect 438 618 454 652
rect 336 568 454 618
rect 336 534 404 568
rect 438 534 454 568
rect 336 485 454 534
rect 336 451 404 485
rect 438 451 454 485
rect 336 435 454 451
rect 248 322 359 356
rect 313 274 359 322
rect 18 258 204 274
rect 18 224 92 258
rect 126 224 204 258
rect 18 158 204 224
rect 18 124 92 158
rect 126 124 204 158
rect 18 113 204 124
rect 18 79 22 113
rect 56 79 94 113
rect 128 79 166 113
rect 200 79 204 113
rect 240 258 359 274
rect 240 224 248 258
rect 282 224 359 258
rect 240 158 359 224
rect 240 124 248 158
rect 282 124 359 158
rect 240 108 359 124
rect 396 258 462 274
rect 396 224 404 258
rect 438 224 462 258
rect 396 158 462 224
rect 396 124 404 158
rect 438 124 462 158
rect 396 113 462 124
rect 18 73 204 79
rect 396 79 402 113
rect 436 79 462 113
rect 396 73 462 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 28 701 62 735
rect 100 701 126 735
rect 126 701 134 735
rect 172 701 206 735
rect 342 701 376 735
rect 414 701 438 735
rect 438 701 448 735
rect 22 79 56 113
rect 94 79 128 113
rect 166 79 200 113
rect 402 79 436 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 831 480 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 480 831
rect 0 791 480 797
rect 0 735 480 763
rect 0 701 28 735
rect 62 701 100 735
rect 134 701 172 735
rect 206 701 342 735
rect 376 701 414 735
rect 448 701 480 735
rect 0 689 480 701
rect 0 113 480 125
rect 0 79 22 113
rect 56 79 94 113
rect 128 79 166 113
rect 200 79 402 113
rect 436 79 480 113
rect 0 51 480 79
rect 0 17 480 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -23 480 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_2
flabel metal1 s 0 51 480 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 0 480 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 689 480 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 480 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 480 814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string LEFsymmetry X Y
string GDS_END 21582
string GDS_START 14604
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016078
<< locali >>
rect 248 961 422 980
rect 248 927 276 961
rect 310 927 360 961
rect 394 927 422 961
rect 248 889 422 927
rect 120 823 186 889
rect 248 855 276 889
rect 310 855 360 889
rect 394 855 422 889
rect 248 841 422 855
rect 484 823 550 889
rect 120 795 160 823
rect 510 795 550 823
rect 41 759 160 795
rect 41 725 60 759
rect 94 725 160 759
rect 41 687 160 725
rect 41 653 60 687
rect 94 653 160 687
rect 41 615 160 653
rect 41 581 60 615
rect 94 581 160 615
rect 41 543 160 581
rect 41 509 60 543
rect 94 509 160 543
rect 41 471 160 509
rect 41 437 60 471
rect 94 437 160 471
rect 41 399 160 437
rect 41 365 60 399
rect 94 365 160 399
rect 41 327 160 365
rect 41 293 60 327
rect 94 293 160 327
rect 41 255 160 293
rect 41 221 60 255
rect 94 221 160 255
rect 41 185 160 221
rect 510 759 629 795
rect 510 725 576 759
rect 610 725 629 759
rect 510 687 629 725
rect 510 653 576 687
rect 610 653 629 687
rect 510 615 629 653
rect 510 581 576 615
rect 610 581 629 615
rect 510 543 629 581
rect 510 509 576 543
rect 610 509 629 543
rect 510 471 629 509
rect 510 437 576 471
rect 610 437 629 471
rect 510 399 629 437
rect 510 365 576 399
rect 610 365 629 399
rect 510 327 629 365
rect 510 293 576 327
rect 610 293 629 327
rect 510 255 629 293
rect 510 221 576 255
rect 610 221 629 255
rect 510 185 629 221
rect 120 157 160 185
rect 510 157 550 185
rect 120 91 186 157
rect 248 125 422 139
rect 248 91 276 125
rect 310 91 360 125
rect 394 91 422 125
rect 484 91 550 157
rect 248 53 422 91
rect 248 19 276 53
rect 310 19 360 53
rect 394 19 422 53
rect 248 0 422 19
<< viali >>
rect 276 927 310 961
rect 360 927 394 961
rect 276 855 310 889
rect 360 855 394 889
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 576 725 610 759
rect 576 653 610 687
rect 576 581 610 615
rect 576 509 610 543
rect 576 437 610 471
rect 576 365 610 399
rect 576 293 610 327
rect 576 221 610 255
rect 276 91 310 125
rect 360 91 394 125
rect 276 19 310 53
rect 360 19 394 53
<< obsli1 >>
rect 212 185 246 795
rect 318 185 352 795
rect 424 185 458 795
<< metal1 >>
rect 250 961 420 980
rect 250 927 276 961
rect 310 927 360 961
rect 394 927 420 961
rect 250 889 420 927
rect 250 855 276 889
rect 310 855 360 889
rect 394 855 420 889
rect 250 843 420 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 570 759 629 771
rect 570 725 576 759
rect 610 725 629 759
rect 570 687 629 725
rect 570 653 576 687
rect 610 653 629 687
rect 570 615 629 653
rect 570 581 576 615
rect 610 581 629 615
rect 570 543 629 581
rect 570 509 576 543
rect 610 509 629 543
rect 570 471 629 509
rect 570 437 576 471
rect 610 437 629 471
rect 570 399 629 437
rect 570 365 576 399
rect 610 365 629 399
rect 570 327 629 365
rect 570 293 576 327
rect 610 293 629 327
rect 570 255 629 293
rect 570 221 576 255
rect 610 221 629 255
rect 570 209 629 221
rect 250 125 420 137
rect 250 91 276 125
rect 310 91 360 125
rect 394 91 420 125
rect 250 53 420 91
rect 250 19 276 53
rect 310 19 360 53
rect 394 19 420 53
rect 250 0 420 19
<< obsm1 >>
rect 203 209 255 771
rect 309 209 361 771
rect 415 209 467 771
<< metal2 >>
rect 14 515 656 771
rect 14 209 656 465
<< labels >>
rlabel viali s 576 725 610 759 6 BULK
port 1 nsew
rlabel viali s 576 653 610 687 6 BULK
port 1 nsew
rlabel viali s 576 581 610 615 6 BULK
port 1 nsew
rlabel viali s 576 509 610 543 6 BULK
port 1 nsew
rlabel viali s 576 437 610 471 6 BULK
port 1 nsew
rlabel viali s 576 365 610 399 6 BULK
port 1 nsew
rlabel viali s 576 293 610 327 6 BULK
port 1 nsew
rlabel viali s 576 221 610 255 6 BULK
port 1 nsew
rlabel viali s 60 725 94 759 6 BULK
port 1 nsew
rlabel viali s 60 653 94 687 6 BULK
port 1 nsew
rlabel viali s 60 581 94 615 6 BULK
port 1 nsew
rlabel viali s 60 509 94 543 6 BULK
port 1 nsew
rlabel viali s 60 437 94 471 6 BULK
port 1 nsew
rlabel viali s 60 365 94 399 6 BULK
port 1 nsew
rlabel viali s 60 293 94 327 6 BULK
port 1 nsew
rlabel viali s 60 221 94 255 6 BULK
port 1 nsew
rlabel locali s 510 795 550 823 6 BULK
port 1 nsew
rlabel locali s 510 185 629 795 6 BULK
port 1 nsew
rlabel locali s 510 157 550 185 6 BULK
port 1 nsew
rlabel locali s 484 823 550 889 6 BULK
port 1 nsew
rlabel locali s 484 91 550 157 6 BULK
port 1 nsew
rlabel locali s 120 823 186 889 6 BULK
port 1 nsew
rlabel locali s 120 795 160 823 6 BULK
port 1 nsew
rlabel locali s 120 157 160 185 6 BULK
port 1 nsew
rlabel locali s 120 91 186 157 6 BULK
port 1 nsew
rlabel locali s 41 185 160 795 6 BULK
port 1 nsew
rlabel metal1 s 570 209 629 771 6 BULK
port 1 nsew
rlabel metal1 s 41 209 100 771 6 BULK
port 1 nsew
rlabel metal2 s 14 515 656 771 6 DRAIN
port 2 nsew
rlabel viali s 360 927 394 961 6 GATE
port 3 nsew
rlabel viali s 360 855 394 889 6 GATE
port 3 nsew
rlabel viali s 360 91 394 125 6 GATE
port 3 nsew
rlabel viali s 360 19 394 53 6 GATE
port 3 nsew
rlabel viali s 276 927 310 961 6 GATE
port 3 nsew
rlabel viali s 276 855 310 889 6 GATE
port 3 nsew
rlabel viali s 276 91 310 125 6 GATE
port 3 nsew
rlabel viali s 276 19 310 53 6 GATE
port 3 nsew
rlabel locali s 248 841 422 980 6 GATE
port 3 nsew
rlabel locali s 248 0 422 139 6 GATE
port 3 nsew
rlabel metal1 s 250 843 420 980 6 GATE
port 3 nsew
rlabel metal1 s 250 0 420 137 6 GATE
port 3 nsew
rlabel metal2 s 14 209 656 465 6 SOURCE
port 4 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 670 980
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9627330
string GDS_START 9612750
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1288 -1260 11168 1731
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_1
timestamp 1633016201
transform 1 0 9880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_0
timestamp 1633016201
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_4
timestamp 1633016201
transform 1 0 8224 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_3
timestamp 1633016201
transform 1 0 6568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_2
timestamp 1633016201
transform 1 0 4912 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_1
timestamp 1633016201
transform 1 0 3256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_0
timestamp 1633016201
transform 1 0 1600 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 9908 471 9908 471 0 FreeSans 300 0 0 0 S
flabel comment s 8252 471 8252 471 0 FreeSans 300 0 0 0 D
flabel comment s 6596 471 6596 471 0 FreeSans 300 0 0 0 S
flabel comment s 4940 471 4940 471 0 FreeSans 300 0 0 0 D
flabel comment s 3284 471 3284 471 0 FreeSans 300 0 0 0 S
flabel comment s 1628 471 1628 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 15441160
string GDS_START 15437708
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016201
<< checkpaint >>
rect -1288 -1260 1448 1731
use sky130_fd_pr__dfl1sd__example_55959141808517  sky130_fd_pr__dfl1sd__example_55959141808517_0
timestamp 1633016201
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808517  sky130_fd_pr__dfl1sd__example_55959141808517_1
timestamp 1633016201
transform 1 0 160 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 188 471 188 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_END 5761016
string GDS_START 5760094
<< end >>

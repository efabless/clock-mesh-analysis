
VVDD      vpwr_0 0  ${VDDD}
VNB       VNB  0  0
VVGND     VGND 0  0

RP_R_0 vpwr_0 vpwr_R_branch_0   ${R_R_BASE}
RP_R_1 vpwr_0 vpwr_R_branch_1   ${R_R_BASE}
RP_R_2 vpwr_0 vpwr_R_branch_2   ${R_R_BASE}
RP_R_3 vpwr_0 vpwr_R_branch_3   ${R_R_BASE}
RP_R_4 vpwr_0 vpwr_R_branch_4   ${R_R_BASE}
RP_R_5 vpwr_0 vpwr_R_branch_5   ${R_R_BASE}
RP_R_6 vpwr_0 vpwr_R_branch_6   ${R_R_BASE}
RP_R_LOAD_0  vpwr_R_branch_0 vpwr_R_0 ${R_R_BUFF}
RP_R_LOAD_1  vpwr_R_branch_1 vpwr_R_1 ${R_R_BUFF}
RP_R_LOAD_2  vpwr_R_branch_2 vpwr_R_2 ${R_R_BUFF}
RP_R_LOAD_3  vpwr_R_branch_3 vpwr_R_3 ${R_R_BUFF}
RP_R_LOAD_4  vpwr_R_branch_4 vpwr_R_4 ${R_R_BUFF}
RP_R_LOAD_5  vpwr_R_branch_5 vpwr_R_5 ${R_R_BUFF}
RP_R_LOAD_6  vpwr_R_branch_6 vpwr_R_6 ${R_R_BUFF}
RP_R_LOAD_7  vpwr_R_branch_0 vpwr_R_7 ${R_R_BUFF}
RP_R_LOAD_8  vpwr_R_branch_1 vpwr_R_8 ${R_R_BUFF}
RP_R_LOAD_9  vpwr_R_branch_2 vpwr_R_9 ${R_R_BUFF}
RP_R_LOAD_10 vpwr_R_branch_3 vpwr_R_10 ${R_R_BUFF}
RP_R_LOAD_11 vpwr_R_branch_4 vpwr_R_11 ${R_R_BUFF}
RP_R_LOAD_12 vpwr_R_branch_5 vpwr_R_12 ${R_R_BUFF}
RP_R_LOAD_13 vpwr_R_branch_6 vpwr_R_13 ${R_R_BUFF}
RP_R_LOAD_14 vpwr_R_branch_0 vpwr_R_14 ${R_R_BUFF}
RP_R_LOAD_15 vpwr_R_branch_1 vpwr_R_15 ${R_R_BUFF}
RP_R_LOAD_16 vpwr_R_branch_2 vpwr_R_16 ${R_R_BUFF}
RP_R_LOAD_17 vpwr_R_branch_3 vpwr_R_17 ${R_R_BUFF}
RP_R_LOAD_18 vpwr_R_branch_4 vpwr_R_18 ${R_R_BUFF}
RP_R_LOAD_19 vpwr_R_branch_5 vpwr_R_19 ${R_R_BUFF}
RP_R_LOAD_20 vpwr_R_branch_6 vpwr_R_20 ${R_R_BUFF}
RP_R_LOAD_21 vpwr_R_branch_0 vpwr_R_21 ${R_R_BUFF}
RP_R_LOAD_22 vpwr_R_branch_1 vpwr_R_22 ${R_R_BUFF}
RP_R_LOAD_23 vpwr_R_branch_2 vpwr_R_23 ${R_R_BUFF}
RP_R_LOAD_24 vpwr_R_branch_3 vpwr_R_24 ${R_R_BUFF}
RP_R_LOAD_25 vpwr_R_branch_4 vpwr_R_25 ${R_R_BUFF}
RP_R_LOAD_26 vpwr_R_branch_5 vpwr_R_26 ${R_R_BUFF}
RP_R_LOAD_27 vpwr_R_branch_6 vpwr_R_27 ${R_R_BUFF}
RP_R_LOAD_28 vpwr_R_branch_0 vpwr_R_28 ${R_R_BUFF}
RP_R_LOAD_29 vpwr_R_branch_1 vpwr_R_29 ${R_R_BUFF}
RP_R_LOAD_30 vpwr_R_branch_2 vpwr_R_30 ${R_R_BUFF}
RP_R_LOAD_31 vpwr_R_branch_3 vpwr_R_31 ${R_R_BUFF}
RP_R_LOAD_32 vpwr_R_branch_4 vpwr_R_32 ${R_R_BUFF}
RP_R_LOAD_33 vpwr_R_branch_5 vpwr_R_33 ${R_R_BUFF}
RP_R_LOAD_34 vpwr_R_branch_6 vpwr_R_34 ${R_R_BUFF}
RP_R_LOAD_35 vpwr_R_branch_0 vpwr_R_35 ${R_R_BUFF}
RP_R_LOAD_36 vpwr_R_branch_1 vpwr_R_36 ${R_R_BUFF}
RP_R_LOAD_37 vpwr_R_branch_2 vpwr_R_37 ${R_R_BUFF}
RP_R_LOAD_38 vpwr_R_branch_3 vpwr_R_38 ${R_R_BUFF}
RP_R_LOAD_39 vpwr_R_branch_4 vpwr_R_39 ${R_R_BUFF}
RP_R_LOAD_40 vpwr_R_branch_5 vpwr_R_40 ${R_R_BUFF}
RP_R_LOAD_41 vpwr_R_branch_6 vpwr_R_41 ${R_R_BUFF}
RP_R_LOAD_42 vpwr_R_branch_0 vpwr_R_42 ${R_R_BUFF}
RP_R_LOAD_43 vpwr_R_branch_1 vpwr_R_43 ${R_R_BUFF}
RP_R_LOAD_44 vpwr_R_branch_2 vpwr_R_44 ${R_R_BUFF}
RP_R_LOAD_45 vpwr_R_branch_3 vpwr_R_45 ${R_R_BUFF}
RP_R_LOAD_46 vpwr_R_branch_4 vpwr_R_46 ${R_R_BUFF}
RP_R_LOAD_47 vpwr_R_branch_5 vpwr_R_47 ${R_R_BUFF}
RP_R_LOAD_48 vpwr_R_branch_6 vpwr_R_48 ${R_R_BUFF}
RP_R_LOAD_49 vpwr_R_branch_0 vpwr_R_49 ${R_R_BUFF}
RP_R_LOAD_50 vpwr_R_branch_1 vpwr_R_50 ${R_R_BUFF}
RP_R_LOAD_51 vpwr_R_branch_2 vpwr_R_51 ${R_R_BUFF}
RP_R_LOAD_52 vpwr_R_branch_3 vpwr_R_52 ${R_R_BUFF}
RP_R_LOAD_53 vpwr_R_branch_4 vpwr_R_53 ${R_R_BUFF}
RP_R_LOAD_54 vpwr_R_branch_5 vpwr_R_54 ${R_R_BUFF}
RP_R_LOAD_55 vpwr_R_branch_6 vpwr_R_55 ${R_R_BUFF}
RP_R_LOAD_56 vpwr_R_branch_0 vpwr_R_56 ${R_R_BUFF}
RP_R_LOAD_57 vpwr_R_branch_1 vpwr_R_57 ${R_R_BUFF}
RP_R_LOAD_58 vpwr_R_branch_2 vpwr_R_58 ${R_R_BUFF}
RP_R_LOAD_59 vpwr_R_branch_3 vpwr_R_59 ${R_R_BUFF}
RP_R_LOAD_60 vpwr_R_branch_4 vpwr_R_60 ${R_R_BUFF}
RP_R_LOAD_61 vpwr_R_branch_5 vpwr_R_61 ${R_R_BUFF}
RP_R_LOAD_62 vpwr_R_branch_6 vpwr_R_62 ${R_R_BUFF}
RP_R_LOAD_63 vpwr_R_branch_0 vpwr_R_63 ${R_R_BUFF}
RP_R_LOAD_64 vpwr_R_branch_1 vpwr_R_64 ${R_R_BUFF}
RP_R_LOAD_65 vpwr_R_branch_2 vpwr_R_65 ${R_R_BUFF}
RP_R_LOAD_66 vpwr_R_branch_3 vpwr_R_66 ${R_R_BUFF}
RP_R_LOAD_67 vpwr_R_branch_4 vpwr_R_67 ${R_R_BUFF}
RP_R_LOAD_68 vpwr_R_branch_5 vpwr_R_68 ${R_R_BUFF}
RP_R_LOAD_69 vpwr_R_branch_6 vpwr_R_69 ${R_R_BUFF}
RP_R_LOAD_70 vpwr_R_branch_0 vpwr_R_70 ${R_R_BUFF}
RP_R_LOAD_71 vpwr_R_branch_1 vpwr_R_71 ${R_R_BUFF}
RP_R_LOAD_72 vpwr_R_branch_2 vpwr_R_72 ${R_R_BUFF}
RP_R_LOAD_73 vpwr_R_branch_3 vpwr_R_73 ${R_R_BUFF}
RP_R_LOAD_74 vpwr_R_branch_4 vpwr_R_74 ${R_R_BUFF}
RP_R_LOAD_75 vpwr_R_branch_5 vpwr_R_75 ${R_R_BUFF}
RP_R_LOAD_76 vpwr_R_branch_6 vpwr_R_76 ${R_R_BUFF}
RP_R_LOAD_77 vpwr_R_branch_0 vpwr_R_77 ${R_R_BUFF}
RP_R_LOAD_78 vpwr_R_branch_1 vpwr_R_78 ${R_R_BUFF}
RP_R_LOAD_79 vpwr_R_branch_2 vpwr_R_79 ${R_R_BUFF}
RP_R_LOAD_80 vpwr_R_branch_3 vpwr_R_80 ${R_R_BUFF}
RP_R_LOAD_81 vpwr_R_branch_4 vpwr_R_81 ${R_R_BUFF}
RP_R_LOAD_82 vpwr_R_branch_5 vpwr_R_82 ${R_R_BUFF}
RP_R_LOAD_83 vpwr_R_branch_6 vpwr_R_83 ${R_R_BUFF}
RP_R_LOAD_84 vpwr_R_branch_0 vpwr_R_84 ${R_R_BUFF}
RP_R_LOAD_85 vpwr_R_branch_1 vpwr_R_85 ${R_R_BUFF}
RP_R_LOAD_86 vpwr_R_branch_2 vpwr_R_86 ${R_R_BUFF}
RP_R_LOAD_87 vpwr_R_branch_3 vpwr_R_87 ${R_R_BUFF}
RP_R_LOAD_88 vpwr_R_branch_4 vpwr_R_88 ${R_R_BUFF}
RP_R_LOAD_89 vpwr_R_branch_5 vpwr_R_89 ${R_R_BUFF}
RP_R_LOAD_90 vpwr_R_branch_6 vpwr_R_90 ${R_R_BUFF}
RP_R_LOAD_91 vpwr_R_branch_0 vpwr_R_91 ${R_R_BUFF}
RP_R_LOAD_92 vpwr_R_branch_1 vpwr_R_92 ${R_R_BUFF}
RP_R_LOAD_93 vpwr_R_branch_2 vpwr_R_93 ${R_R_BUFF}
RP_R_LOAD_94 vpwr_R_branch_3 vpwr_R_94 ${R_R_BUFF}
RP_R_LOAD_95 vpwr_R_branch_4 vpwr_R_95 ${R_R_BUFF}
RP_R_LOAD_96 vpwr_R_branch_5 vpwr_R_96 ${R_R_BUFF}
RP_R_LOAD_97 vpwr_R_branch_6 vpwr_R_97 ${R_R_BUFF}
RP_R_LOAD_98 vpwr_R_branch_0 vpwr_R_98 ${R_R_BUFF}
RP_R_LOAD_99 vpwr_R_branch_1 vpwr_R_99 ${R_R_BUFF}
RP_R_LOAD_100 vpwr_R_branch_2 vpwr_R_100 ${R_R_BUFF}
RP_R_LOAD_101 vpwr_R_branch_3 vpwr_R_101 ${R_R_BUFF}
RP_R_LOAD_102 vpwr_R_branch_4 vpwr_R_102 ${R_R_BUFF}
RP_R_LOAD_103 vpwr_R_branch_5 vpwr_R_103 ${R_R_BUFF}
RP_R_LOAD_104 vpwr_R_branch_6 vpwr_R_104 ${R_R_BUFF}
RP_R_LOAD_105 vpwr_R_branch_0 vpwr_R_105 ${R_R_BUFF}
RP_R_LOAD_106 vpwr_R_branch_1 vpwr_R_106 ${R_R_BUFF}
RP_R_LOAD_107 vpwr_R_branch_2 vpwr_R_107 ${R_R_BUFF}
RP_R_LOAD_108 vpwr_R_branch_3 vpwr_R_108 ${R_R_BUFF}
RP_R_LOAD_109 vpwr_R_branch_4 vpwr_R_109 ${R_R_BUFF}
RP_R_LOAD_110 vpwr_R_branch_5 vpwr_R_110 ${R_R_BUFF}
RP_R_LOAD_111 vpwr_R_branch_6 vpwr_R_111 ${R_R_BUFF}
RP_R_LOAD_112 vpwr_R_branch_0 vpwr_R_112 ${R_R_BUFF}
RP_R_LOAD_113 vpwr_R_branch_1 vpwr_R_113 ${R_R_BUFF}
RP_R_LOAD_114 vpwr_R_branch_2 vpwr_R_114 ${R_R_BUFF}
RP_R_LOAD_115 vpwr_R_branch_3 vpwr_R_115 ${R_R_BUFF}
RP_R_LOAD_116 vpwr_R_branch_4 vpwr_R_116 ${R_R_BUFF}
RP_R_LOAD_117 vpwr_R_branch_5 vpwr_R_117 ${R_R_BUFF}
RP_R_LOAD_118 vpwr_R_branch_6 vpwr_R_118 ${R_R_BUFF}
RP_R_LOAD_119 vpwr_R_branch_0 vpwr_R_119 ${R_R_BUFF}
RP_R_LOAD_120 vpwr_R_branch_1 vpwr_R_120 ${R_R_BUFF}
RP_R_LOAD_121 vpwr_R_branch_2 vpwr_R_121 ${R_R_BUFF}
RP_R_LOAD_122 vpwr_R_branch_3 vpwr_R_122 ${R_R_BUFF}
RP_R_LOAD_123 vpwr_R_branch_4 vpwr_R_123 ${R_R_BUFF}
RP_R_LOAD_124 vpwr_R_branch_5 vpwr_R_124 ${R_R_BUFF}
RP_R_LOAD_125 vpwr_R_branch_6 vpwr_R_125 ${R_R_BUFF}
RP_R_LOAD_126 vpwr_R_branch_0 vpwr_R_126 ${R_R_BUFF}
RP_R_LOAD_127 vpwr_R_branch_1 vpwr_R_127 ${R_R_BUFF}
RP_R_LOAD_128 vpwr_R_branch_2 vpwr_R_128 ${R_R_BUFF}
RP_R_LOAD_129 vpwr_R_branch_3 vpwr_R_129 ${R_R_BUFF}
RP_R_LOAD_130 vpwr_R_branch_4 vpwr_R_130 ${R_R_BUFF}
RP_R_LOAD_131 vpwr_R_branch_5 vpwr_R_131 ${R_R_BUFF}
RP_R_LOAD_132 vpwr_R_branch_6 vpwr_R_132 ${R_R_BUFF}
RP_R_LOAD_133 vpwr_R_branch_0 vpwr_R_133 ${R_R_BUFF}
RP_R_LOAD_134 vpwr_R_branch_1 vpwr_R_134 ${R_R_BUFF}
RP_R_LOAD_135 vpwr_R_branch_2 vpwr_R_135 ${R_R_BUFF}
RP_R_LOAD_136 vpwr_R_branch_3 vpwr_R_136 ${R_R_BUFF}
RP_R_LOAD_137 vpwr_R_branch_4 vpwr_R_137 ${R_R_BUFF}
RP_R_LOAD_138 vpwr_R_branch_5 vpwr_R_138 ${R_R_BUFF}
RP_R_LOAD_139 vpwr_R_branch_6 vpwr_R_139 ${R_R_BUFF}
RP_R_LOAD_140 vpwr_R_branch_0 vpwr_R_140 ${R_R_BUFF}
RP_R_LOAD_141 vpwr_R_branch_1 vpwr_R_141 ${R_R_BUFF}
RP_R_LOAD_142 vpwr_R_branch_2 vpwr_R_142 ${R_R_BUFF}
RP_R_LOAD_143 vpwr_R_branch_3 vpwr_R_143 ${R_R_BUFF}
RP_R_LOAD_144 vpwr_R_branch_4 vpwr_R_144 ${R_R_BUFF}
RP_R_LOAD_145 vpwr_R_branch_5 vpwr_R_145 ${R_R_BUFF}
RP_R_LOAD_146 vpwr_R_branch_6 vpwr_R_146 ${R_R_BUFF}
RP_R_LOAD_147 vpwr_R_branch_0 vpwr_R_147 ${R_R_BUFF}
RP_R_LOAD_148 vpwr_R_branch_1 vpwr_R_148 ${R_R_BUFF}
RP_R_LOAD_149 vpwr_R_branch_2 vpwr_R_149 ${R_R_BUFF}
RP_R_LOAD_150 vpwr_R_branch_3 vpwr_R_150 ${R_R_BUFF}
RP_R_LOAD_151 vpwr_R_branch_4 vpwr_R_151 ${R_R_BUFF}
RP_R_LOAD_152 vpwr_R_branch_5 vpwr_R_152 ${R_R_BUFF}
RP_R_LOAD_153 vpwr_R_branch_6 vpwr_R_153 ${R_R_BUFF}
RP_R_LOAD_154 vpwr_R_branch_0 vpwr_R_154 ${R_R_BUFF}
RP_R_LOAD_155 vpwr_R_branch_1 vpwr_R_155 ${R_R_BUFF}
RP_R_LOAD_156 vpwr_R_branch_2 vpwr_R_156 ${R_R_BUFF}
RP_R_LOAD_157 vpwr_R_branch_3 vpwr_R_157 ${R_R_BUFF}
RP_R_LOAD_158 vpwr_R_branch_4 vpwr_R_158 ${R_R_BUFF}
RP_R_LOAD_159 vpwr_R_branch_5 vpwr_R_159 ${R_R_BUFF}
RP_R_LOAD_160 vpwr_R_branch_6 vpwr_R_160 ${R_R_BUFF}
RP_R_LOAD_161 vpwr_R_branch_0 vpwr_R_161 ${R_R_BUFF}
RP_R_LOAD_162 vpwr_R_branch_1 vpwr_R_162 ${R_R_BUFF}
RP_R_LOAD_163 vpwr_R_branch_2 vpwr_R_163 ${R_R_BUFF}
RP_R_LOAD_164 vpwr_R_branch_3 vpwr_R_164 ${R_R_BUFF}
RP_R_LOAD_165 vpwr_R_branch_4 vpwr_R_165 ${R_R_BUFF}
RP_R_LOAD_166 vpwr_R_branch_5 vpwr_R_166 ${R_R_BUFF}
RP_R_LOAD_167 vpwr_R_branch_6 vpwr_R_167 ${R_R_BUFF}
RP_R_LOAD_168 vpwr_R_branch_0 vpwr_R_168 ${R_R_BUFF}
RP_R_LOAD_169 vpwr_R_branch_1 vpwr_R_169 ${R_R_BUFF}
RP_R_LOAD_170 vpwr_R_branch_2 vpwr_R_170 ${R_R_BUFF}
RP_R_LOAD_171 vpwr_R_branch_3 vpwr_R_171 ${R_R_BUFF}
RP_R_LOAD_172 vpwr_R_branch_4 vpwr_R_172 ${R_R_BUFF}
RP_R_LOAD_173 vpwr_R_branch_5 vpwr_R_173 ${R_R_BUFF}
RP_R_LOAD_174 vpwr_R_branch_6 vpwr_R_174 ${R_R_BUFF}
RP_R_LOAD_175 vpwr_R_branch_0 vpwr_R_175 ${R_R_BUFF}
RP_R_LOAD_176 vpwr_R_branch_1 vpwr_R_176 ${R_R_BUFF}
RP_R_LOAD_177 vpwr_R_branch_2 vpwr_R_177 ${R_R_BUFF}
RP_R_LOAD_178 vpwr_R_branch_3 vpwr_R_178 ${R_R_BUFF}
RP_R_LOAD_179 vpwr_R_branch_4 vpwr_R_179 ${R_R_BUFF}
RP_R_LOAD_180 vpwr_R_branch_5 vpwr_R_180 ${R_R_BUFF}
RP_R_LOAD_181 vpwr_R_branch_6 vpwr_R_181 ${R_R_BUFF}
RP_R_LOAD_182 vpwr_R_branch_0 vpwr_R_182 ${R_R_BUFF}
RP_R_LOAD_183 vpwr_R_branch_1 vpwr_R_183 ${R_R_BUFF}
RP_R_LOAD_184 vpwr_R_branch_2 vpwr_R_184 ${R_R_BUFF}
RP_R_LOAD_185 vpwr_R_branch_3 vpwr_R_185 ${R_R_BUFF}
RP_R_LOAD_186 vpwr_R_branch_4 vpwr_R_186 ${R_R_BUFF}
RP_R_LOAD_187 vpwr_R_branch_5 vpwr_R_187 ${R_R_BUFF}
RP_R_LOAD_188 vpwr_R_branch_6 vpwr_R_188 ${R_R_BUFF}
RP_R_LOAD_189 vpwr_R_branch_0 vpwr_R_189 ${R_R_BUFF}
RP_R_LOAD_190 vpwr_R_branch_1 vpwr_R_190 ${R_R_BUFF}
RP_R_LOAD_191 vpwr_R_branch_2 vpwr_R_191 ${R_R_BUFF}
RP_R_LOAD_192 vpwr_R_branch_3 vpwr_R_192 ${R_R_BUFF}
RP_R_LOAD_193 vpwr_R_branch_4 vpwr_R_193 ${R_R_BUFF}
RP_R_LOAD_194 vpwr_R_branch_5 vpwr_R_194 ${R_R_BUFF}
RP_R_LOAD_195 vpwr_R_branch_6 vpwr_R_195 ${R_R_BUFF}
RP_R_LOAD_196 vpwr_R_branch_0 vpwr_R_196 ${R_R_BUFF}
RP_R_LOAD_197 vpwr_R_branch_1 vpwr_R_197 ${R_R_BUFF}
RP_R_LOAD_198 vpwr_R_branch_2 vpwr_R_198 ${R_R_BUFF}
RP_R_LOAD_199 vpwr_R_branch_3 vpwr_R_199 ${R_R_BUFF}
RP_R_LOAD_200 vpwr_R_branch_4 vpwr_R_200 ${R_R_BUFF}
RP_R_LOAD_201 vpwr_R_branch_5 vpwr_R_201 ${R_R_BUFF}
RP_R_LOAD_202 vpwr_R_branch_6 vpwr_R_202 ${R_R_BUFF}
RP_R_LOAD_203 vpwr_R_branch_0 vpwr_R_203 ${R_R_BUFF}
RP_R_LOAD_204 vpwr_R_branch_1 vpwr_R_204 ${R_R_BUFF}
RP_R_LOAD_205 vpwr_R_branch_2 vpwr_R_205 ${R_R_BUFF}
RP_R_LOAD_206 vpwr_R_branch_3 vpwr_R_206 ${R_R_BUFF}
RP_R_LOAD_207 vpwr_R_branch_4 vpwr_R_207 ${R_R_BUFF}
RP_R_LOAD_208 vpwr_R_branch_5 vpwr_R_208 ${R_R_BUFF}
RP_R_LOAD_209 vpwr_R_branch_6 vpwr_R_209 ${R_R_BUFF}
RP_R_LOAD_210 vpwr_R_branch_0 vpwr_R_210 ${R_R_BUFF}
RP_R_LOAD_211 vpwr_R_branch_1 vpwr_R_211 ${R_R_BUFF}
RP_R_LOAD_212 vpwr_R_branch_2 vpwr_R_212 ${R_R_BUFF}
RP_R_LOAD_213 vpwr_R_branch_3 vpwr_R_213 ${R_R_BUFF}
RP_R_LOAD_214 vpwr_R_branch_4 vpwr_R_214 ${R_R_BUFF}
RP_R_LOAD_215 vpwr_R_branch_5 vpwr_R_215 ${R_R_BUFF}
RP_R_LOAD_216 vpwr_R_branch_6 vpwr_R_216 ${R_R_BUFF}
RP_R_LOAD_217 vpwr_R_branch_0 vpwr_R_217 ${R_R_BUFF}
RP_R_LOAD_218 vpwr_R_branch_1 vpwr_R_218 ${R_R_BUFF}
RP_R_LOAD_219 vpwr_R_branch_2 vpwr_R_219 ${R_R_BUFF}
RP_R_LOAD_220 vpwr_R_branch_3 vpwr_R_220 ${R_R_BUFF}
RP_R_LOAD_221 vpwr_R_branch_4 vpwr_R_221 ${R_R_BUFF}
RP_R_LOAD_222 vpwr_R_branch_5 vpwr_R_222 ${R_R_BUFF}
RP_R_LOAD_223 vpwr_R_branch_6 vpwr_R_223 ${R_R_BUFF}
RP_R_LOAD_224 vpwr_R_branch_0 vpwr_R_224 ${R_R_BUFF}
RP_R_LOAD_225 vpwr_R_branch_1 vpwr_R_225 ${R_R_BUFF}
RP_R_LOAD_226 vpwr_R_branch_2 vpwr_R_226 ${R_R_BUFF}
RP_R_LOAD_227 vpwr_R_branch_3 vpwr_R_227 ${R_R_BUFF}
RP_R_LOAD_228 vpwr_R_branch_4 vpwr_R_228 ${R_R_BUFF}
RP_R_LOAD_229 vpwr_R_branch_5 vpwr_R_229 ${R_R_BUFF}
RP_R_LOAD_230 vpwr_R_branch_6 vpwr_R_230 ${R_R_BUFF}
RP_R_LOAD_231 vpwr_R_branch_0 vpwr_R_231 ${R_R_BUFF}
RP_R_LOAD_232 vpwr_R_branch_1 vpwr_R_232 ${R_R_BUFF}
RP_R_LOAD_233 vpwr_R_branch_2 vpwr_R_233 ${R_R_BUFF}
RP_R_LOAD_234 vpwr_R_branch_3 vpwr_R_234 ${R_R_BUFF}
RP_R_LOAD_235 vpwr_R_branch_4 vpwr_R_235 ${R_R_BUFF}
RP_R_LOAD_236 vpwr_R_branch_5 vpwr_R_236 ${R_R_BUFF}
RP_R_LOAD_237 vpwr_R_branch_6 vpwr_R_237 ${R_R_BUFF}
RP_R_LOAD_238 vpwr_R_branch_0 vpwr_R_238 ${R_R_BUFF}
RP_R_LOAD_239 vpwr_R_branch_1 vpwr_R_239 ${R_R_BUFF}
RP_R_LOAD_240 vpwr_R_branch_2 vpwr_R_240 ${R_R_BUFF}
RP_R_LOAD_241 vpwr_R_branch_3 vpwr_R_241 ${R_R_BUFF}
RP_R_LOAD_242 vpwr_R_branch_4 vpwr_R_242 ${R_R_BUFF}
RP_R_LOAD_243 vpwr_R_branch_5 vpwr_R_243 ${R_R_BUFF}
RP_R_LOAD_244 vpwr_R_branch_6 vpwr_R_244 ${R_R_BUFF}
RP_R_LOAD_245 vpwr_R_branch_0 vpwr_R_245 ${R_R_BUFF}
RP_R_LOAD_246 vpwr_R_branch_1 vpwr_R_246 ${R_R_BUFF}
RP_R_LOAD_247 vpwr_R_branch_2 vpwr_R_247 ${R_R_BUFF}
RP_R_LOAD_248 vpwr_R_branch_3 vpwr_R_248 ${R_R_BUFF}
RP_R_LOAD_249 vpwr_R_branch_4 vpwr_R_249 ${R_R_BUFF}
RP_R_LOAD_250 vpwr_R_branch_5 vpwr_R_250 ${R_R_BUFF}
RP_R_LOAD_251 vpwr_R_branch_6 vpwr_R_251 ${R_R_BUFF}
RP_R_LOAD_252 vpwr_R_branch_0 vpwr_R_252 ${R_R_BUFF}
RP_R_LOAD_253 vpwr_R_branch_1 vpwr_R_253 ${R_R_BUFF}
RP_R_LOAD_254 vpwr_R_branch_2 vpwr_R_254 ${R_R_BUFF}
RP_R_LOAD_255 vpwr_R_branch_3 vpwr_R_255 ${R_R_BUFF}
RP_R_LOAD_256 vpwr_R_branch_4 vpwr_R_256 ${R_R_BUFF}
RP_R_LOAD_257 vpwr_R_branch_5 vpwr_R_257 ${R_R_BUFF}
RP_R_LOAD_258 vpwr_R_branch_6 vpwr_R_258 ${R_R_BUFF}
RP_R_LOAD_259 vpwr_R_branch_0 vpwr_R_259 ${R_R_BUFF}
RP_R_LOAD_260 vpwr_R_branch_1 vpwr_R_260 ${R_R_BUFF}
RP_R_LOAD_261 vpwr_R_branch_2 vpwr_R_261 ${R_R_BUFF}
RP_R_LOAD_262 vpwr_R_branch_3 vpwr_R_262 ${R_R_BUFF}
RP_R_LOAD_263 vpwr_R_branch_4 vpwr_R_263 ${R_R_BUFF}
RP_R_LOAD_264 vpwr_R_branch_5 vpwr_R_264 ${R_R_BUFF}
RP_R_LOAD_265 vpwr_R_branch_6 vpwr_R_265 ${R_R_BUFF}
RP_R_LOAD_266 vpwr_R_branch_0 vpwr_R_266 ${R_R_BUFF}
RP_R_LOAD_267 vpwr_R_branch_1 vpwr_R_267 ${R_R_BUFF}
RP_R_LOAD_268 vpwr_R_branch_2 vpwr_R_268 ${R_R_BUFF}
RP_R_LOAD_269 vpwr_R_branch_3 vpwr_R_269 ${R_R_BUFF}
RP_R_LOAD_270 vpwr_R_branch_4 vpwr_R_270 ${R_R_BUFF}
RP_R_LOAD_271 vpwr_R_branch_5 vpwr_R_271 ${R_R_BUFF}
RP_R_LOAD_272 vpwr_R_branch_6 vpwr_R_272 ${R_R_BUFF}
RP_R_LOAD_273 vpwr_R_branch_0 vpwr_R_273 ${R_R_BUFF}
RP_R_LOAD_274 vpwr_R_branch_1 vpwr_R_274 ${R_R_BUFF}
RP_R_LOAD_275 vpwr_R_branch_2 vpwr_R_275 ${R_R_BUFF}
RP_R_LOAD_276 vpwr_R_branch_3 vpwr_R_276 ${R_R_BUFF}
RP_R_LOAD_277 vpwr_R_branch_4 vpwr_R_277 ${R_R_BUFF}
RP_R_LOAD_278 vpwr_R_branch_5 vpwr_R_278 ${R_R_BUFF}
RP_R_LOAD_279 vpwr_R_branch_6 vpwr_R_279 ${R_R_BUFF}
RP_R_LOAD_280 vpwr_R_branch_0 vpwr_R_280 ${R_R_BUFF}
RP_R_LOAD_281 vpwr_R_branch_1 vpwr_R_281 ${R_R_BUFF}
RP_R_LOAD_282 vpwr_R_branch_2 vpwr_R_282 ${R_R_BUFF}
RP_R_LOAD_283 vpwr_R_branch_3 vpwr_R_283 ${R_R_BUFF}
RP_R_LOAD_284 vpwr_R_branch_4 vpwr_R_284 ${R_R_BUFF}
RP_R_LOAD_285 vpwr_R_branch_5 vpwr_R_285 ${R_R_BUFF}
RP_R_LOAD_286 vpwr_R_branch_6 vpwr_R_286 ${R_R_BUFF}
RP_R_LOAD_287 vpwr_R_branch_0 vpwr_R_287 ${R_R_BUFF}
RP_R_LOAD_288 vpwr_R_branch_1 vpwr_R_288 ${R_R_BUFF}
RP_R_LOAD_289 vpwr_R_branch_2 vpwr_R_289 ${R_R_BUFF}
RP_R_LOAD_290 vpwr_R_branch_3 vpwr_R_290 ${R_R_BUFF}
RP_R_LOAD_291 vpwr_R_branch_4 vpwr_R_291 ${R_R_BUFF}
RP_R_LOAD_292 vpwr_R_branch_5 vpwr_R_292 ${R_R_BUFF}
RP_R_LOAD_293 vpwr_R_branch_6 vpwr_R_293 ${R_R_BUFF}
RP_R_LOAD_294 vpwr_R_branch_0 vpwr_R_294 ${R_R_BUFF}
RP_R_LOAD_295 vpwr_R_branch_1 vpwr_R_295 ${R_R_BUFF}
RP_R_LOAD_296 vpwr_R_branch_2 vpwr_R_296 ${R_R_BUFF}
RP_R_LOAD_297 vpwr_R_branch_3 vpwr_R_297 ${R_R_BUFF}
RP_R_LOAD_298 vpwr_R_branch_4 vpwr_R_298 ${R_R_BUFF}
RP_R_LOAD_299 vpwr_R_branch_5 vpwr_R_299 ${R_R_BUFF}
RP_R_LOAD_300 vpwr_R_branch_6 vpwr_R_300 ${R_R_BUFF}
RP_R_LOAD_301 vpwr_R_branch_0 vpwr_R_301 ${R_R_BUFF}
RP_R_LOAD_302 vpwr_R_branch_1 vpwr_R_302 ${R_R_BUFF}
RP_R_LOAD_303 vpwr_R_branch_2 vpwr_R_303 ${R_R_BUFF}
RP_R_LOAD_304 vpwr_R_branch_3 vpwr_R_304 ${R_R_BUFF}
RP_R_LOAD_305 vpwr_R_branch_4 vpwr_R_305 ${R_R_BUFF}
RP_R_LOAD_306 vpwr_R_branch_5 vpwr_R_306 ${R_R_BUFF}
RP_R_LOAD_307 vpwr_R_branch_6 vpwr_R_307 ${R_R_BUFF}
RP_R_LOAD_308 vpwr_R_branch_0 vpwr_R_308 ${R_R_BUFF}
RP_R_LOAD_309 vpwr_R_branch_1 vpwr_R_309 ${R_R_BUFF}
RP_R_LOAD_310 vpwr_R_branch_2 vpwr_R_310 ${R_R_BUFF}
RP_R_LOAD_311 vpwr_R_branch_3 vpwr_R_311 ${R_R_BUFF}
RP_R_LOAD_312 vpwr_R_branch_4 vpwr_R_312 ${R_R_BUFF}
RP_R_LOAD_313 vpwr_R_branch_5 vpwr_R_313 ${R_R_BUFF}
RP_R_LOAD_314 vpwr_R_branch_6 vpwr_R_314 ${R_R_BUFF}
RP_R_LOAD_315 vpwr_R_branch_0 vpwr_R_315 ${R_R_BUFF}
RP_R_LOAD_316 vpwr_R_branch_1 vpwr_R_316 ${R_R_BUFF}
RP_R_LOAD_317 vpwr_R_branch_2 vpwr_R_317 ${R_R_BUFF}
RP_R_LOAD_318 vpwr_R_branch_3 vpwr_R_318 ${R_R_BUFF}
RP_R_LOAD_319 vpwr_R_branch_4 vpwr_R_319 ${R_R_BUFF}
RP_R_LOAD_320 vpwr_R_branch_5 vpwr_R_320 ${R_R_BUFF}
RP_R_LOAD_321 vpwr_R_branch_6 vpwr_R_321 ${R_R_BUFF}
RP_R_LOAD_322 vpwr_R_branch_0 vpwr_R_322 ${R_R_BUFF}
RP_R_LOAD_323 vpwr_R_branch_1 vpwr_R_323 ${R_R_BUFF}
RP_R_LOAD_324 vpwr_R_branch_2 vpwr_R_324 ${R_R_BUFF}
RP_R_LOAD_325 vpwr_R_branch_3 vpwr_R_325 ${R_R_BUFF}
RP_R_LOAD_326 vpwr_R_branch_4 vpwr_R_326 ${R_R_BUFF}
RP_R_LOAD_327 vpwr_R_branch_5 vpwr_R_327 ${R_R_BUFF}
RP_R_LOAD_328 vpwr_R_branch_6 vpwr_R_328 ${R_R_BUFF}
RP_R_LOAD_329 vpwr_R_branch_0 vpwr_R_329 ${R_R_BUFF}
RP_R_LOAD_330 vpwr_R_branch_1 vpwr_R_330 ${R_R_BUFF}
RP_R_LOAD_331 vpwr_R_branch_2 vpwr_R_331 ${R_R_BUFF}
RP_R_LOAD_332 vpwr_R_branch_3 vpwr_R_332 ${R_R_BUFF}
RP_R_LOAD_333 vpwr_R_branch_4 vpwr_R_333 ${R_R_BUFF}
RP_R_LOAD_334 vpwr_R_branch_5 vpwr_R_334 ${R_R_BUFF}
RP_R_LOAD_335 vpwr_R_branch_6 vpwr_R_335 ${R_R_BUFF}
RP_R_LOAD_336 vpwr_R_branch_0 vpwr_R_336 ${R_R_BUFF}
RP_R_LOAD_337 vpwr_R_branch_1 vpwr_R_337 ${R_R_BUFF}
RP_R_LOAD_338 vpwr_R_branch_2 vpwr_R_338 ${R_R_BUFF}
RP_R_LOAD_339 vpwr_R_branch_3 vpwr_R_339 ${R_R_BUFF}
RP_R_LOAD_340 vpwr_R_branch_4 vpwr_R_340 ${R_R_BUFF}
RP_R_LOAD_341 vpwr_R_branch_5 vpwr_R_341 ${R_R_BUFF}
RP_R_LOAD_342 vpwr_R_branch_6 vpwr_R_342 ${R_R_BUFF}
RP_R_LOAD_343 vpwr_R_branch_0 vpwr_R_343 ${R_R_BUFF}
RP_R_LOAD_344 vpwr_R_branch_1 vpwr_R_344 ${R_R_BUFF}
RP_R_LOAD_345 vpwr_R_branch_2 vpwr_R_345 ${R_R_BUFF}
RP_R_LOAD_346 vpwr_R_branch_3 vpwr_R_346 ${R_R_BUFF}
RP_R_LOAD_347 vpwr_R_branch_4 vpwr_R_347 ${R_R_BUFF}
RP_R_LOAD_348 vpwr_R_branch_5 vpwr_R_348 ${R_R_BUFF}
RP_R_LOAD_349 vpwr_R_branch_6 vpwr_R_349 ${R_R_BUFF}
RP_R_LOAD_350 vpwr_R_branch_0 vpwr_R_350 ${R_R_BUFF}
RP_R_LOAD_351 vpwr_R_branch_1 vpwr_R_351 ${R_R_BUFF}
RP_R_LOAD_352 vpwr_R_branch_2 vpwr_R_352 ${R_R_BUFF}
RP_R_LOAD_353 vpwr_R_branch_3 vpwr_R_353 ${R_R_BUFF}
RP_R_LOAD_354 vpwr_R_branch_4 vpwr_R_354 ${R_R_BUFF}
RP_R_LOAD_355 vpwr_R_branch_5 vpwr_R_355 ${R_R_BUFF}
RP_R_LOAD_356 vpwr_R_branch_6 vpwr_R_356 ${R_R_BUFF}
RP_R_LOAD_357 vpwr_R_branch_0 vpwr_R_357 ${R_R_BUFF}
RP_R_LOAD_358 vpwr_R_branch_1 vpwr_R_358 ${R_R_BUFF}
RP_R_LOAD_359 vpwr_R_branch_2 vpwr_R_359 ${R_R_BUFF}
RP_R_LOAD_360 vpwr_R_branch_3 vpwr_R_360 ${R_R_BUFF}
RP_R_LOAD_361 vpwr_R_branch_4 vpwr_R_361 ${R_R_BUFF}
RP_R_LOAD_362 vpwr_R_branch_5 vpwr_R_362 ${R_R_BUFF}
RP_R_LOAD_363 vpwr_R_branch_6 vpwr_R_363 ${R_R_BUFF}
RP_R_LOAD_364 vpwr_R_branch_0 vpwr_R_364 ${R_R_BUFF}
RP_R_LOAD_365 vpwr_R_branch_1 vpwr_R_365 ${R_R_BUFF}
RP_R_LOAD_366 vpwr_R_branch_2 vpwr_R_366 ${R_R_BUFF}
RP_R_LOAD_367 vpwr_R_branch_3 vpwr_R_367 ${R_R_BUFF}
RP_R_LOAD_368 vpwr_R_branch_4 vpwr_R_368 ${R_R_BUFF}
RP_R_LOAD_369 vpwr_R_branch_5 vpwr_R_369 ${R_R_BUFF}
RP_R_LOAD_370 vpwr_R_branch_6 vpwr_R_370 ${R_R_BUFF}
RP_R_LOAD_371 vpwr_R_branch_0 vpwr_R_371 ${R_R_BUFF}
RP_R_LOAD_372 vpwr_R_branch_1 vpwr_R_372 ${R_R_BUFF}
RP_R_LOAD_373 vpwr_R_branch_2 vpwr_R_373 ${R_R_BUFF}
RP_R_LOAD_374 vpwr_R_branch_3 vpwr_R_374 ${R_R_BUFF}
RP_R_LOAD_375 vpwr_R_branch_4 vpwr_R_375 ${R_R_BUFF}
RP_R_LOAD_376 vpwr_R_branch_5 vpwr_R_376 ${R_R_BUFF}
RP_R_LOAD_377 vpwr_R_branch_6 vpwr_R_377 ${R_R_BUFF}
RP_R_LOAD_378 vpwr_R_branch_0 vpwr_R_378 ${R_R_BUFF}
RP_R_LOAD_379 vpwr_R_branch_1 vpwr_R_379 ${R_R_BUFF}
RP_R_LOAD_380 vpwr_R_branch_2 vpwr_R_380 ${R_R_BUFF}
RP_R_LOAD_381 vpwr_R_branch_3 vpwr_R_381 ${R_R_BUFF}
RP_R_LOAD_382 vpwr_R_branch_4 vpwr_R_382 ${R_R_BUFF}
RP_R_LOAD_383 vpwr_R_branch_5 vpwr_R_383 ${R_R_BUFF}
RP_R_LOAD_384 vpwr_R_branch_6 vpwr_R_384 ${R_R_BUFF}
RP_R_LOAD_385 vpwr_R_branch_0 vpwr_R_385 ${R_R_BUFF}
RP_R_LOAD_386 vpwr_R_branch_1 vpwr_R_386 ${R_R_BUFF}
RP_R_LOAD_387 vpwr_R_branch_2 vpwr_R_387 ${R_R_BUFF}
RP_R_LOAD_388 vpwr_R_branch_3 vpwr_R_388 ${R_R_BUFF}
RP_R_LOAD_389 vpwr_R_branch_4 vpwr_R_389 ${R_R_BUFF}
RP_R_LOAD_390 vpwr_R_branch_5 vpwr_R_390 ${R_R_BUFF}
RP_R_LOAD_391 vpwr_R_branch_6 vpwr_R_391 ${R_R_BUFF}
RP_R_LOAD_392 vpwr_R_branch_0 vpwr_R_392 ${R_R_BUFF}
RP_R_LOAD_393 vpwr_R_branch_1 vpwr_R_393 ${R_R_BUFF}
RP_R_LOAD_394 vpwr_R_branch_2 vpwr_R_394 ${R_R_BUFF}
RP_R_LOAD_395 vpwr_R_branch_3 vpwr_R_395 ${R_R_BUFF}
RP_R_LOAD_396 vpwr_R_branch_4 vpwr_R_396 ${R_R_BUFF}
RP_R_LOAD_397 vpwr_R_branch_5 vpwr_R_397 ${R_R_BUFF}
RP_R_LOAD_398 vpwr_R_branch_6 vpwr_R_398 ${R_R_BUFF}
RP_R_LOAD_399 vpwr_R_branch_0 vpwr_R_399 ${R_R_BUFF}
RP_R_LOAD_400 vpwr_R_branch_1 vpwr_R_400 ${R_R_BUFF}
RP_R_LOAD_401 vpwr_R_branch_2 vpwr_R_401 ${R_R_BUFF}
RP_R_LOAD_402 vpwr_R_branch_3 vpwr_R_402 ${R_R_BUFF}
RP_R_LOAD_403 vpwr_R_branch_4 vpwr_R_403 ${R_R_BUFF}
RP_R_LOAD_404 vpwr_R_branch_5 vpwr_R_404 ${R_R_BUFF}
RP_R_LOAD_405 vpwr_R_branch_6 vpwr_R_405 ${R_R_BUFF}
RP_R_LOAD_406 vpwr_R_branch_0 vpwr_R_406 ${R_R_BUFF}
RP_R_LOAD_407 vpwr_R_branch_1 vpwr_R_407 ${R_R_BUFF}
RP_R_LOAD_408 vpwr_R_branch_2 vpwr_R_408 ${R_R_BUFF}
RP_R_LOAD_409 vpwr_R_branch_3 vpwr_R_409 ${R_R_BUFF}
RP_R_LOAD_410 vpwr_R_branch_4 vpwr_R_410 ${R_R_BUFF}
RP_R_LOAD_411 vpwr_R_branch_5 vpwr_R_411 ${R_R_BUFF}
RP_R_LOAD_412 vpwr_R_branch_6 vpwr_R_412 ${R_R_BUFF}
RP_R_LOAD_413 vpwr_R_branch_0 vpwr_R_413 ${R_R_BUFF}
RP_R_LOAD_414 vpwr_R_branch_1 vpwr_R_414 ${R_R_BUFF}
RP_R_LOAD_415 vpwr_R_branch_2 vpwr_R_415 ${R_R_BUFF}
RP_R_LOAD_416 vpwr_R_branch_3 vpwr_R_416 ${R_R_BUFF}
RP_R_LOAD_417 vpwr_R_branch_4 vpwr_R_417 ${R_R_BUFF}
RP_R_LOAD_418 vpwr_R_branch_5 vpwr_R_418 ${R_R_BUFF}
RP_R_LOAD_419 vpwr_R_branch_6 vpwr_R_419 ${R_R_BUFF}
RP_R_LOAD_420 vpwr_R_branch_0 vpwr_R_420 ${R_R_BUFF}
RP_R_LOAD_421 vpwr_R_branch_1 vpwr_R_421 ${R_R_BUFF}
RP_R_LOAD_422 vpwr_R_branch_2 vpwr_R_422 ${R_R_BUFF}
RP_R_LOAD_423 vpwr_R_branch_3 vpwr_R_423 ${R_R_BUFF}
RP_R_LOAD_424 vpwr_R_branch_4 vpwr_R_424 ${R_R_BUFF}
RP_R_LOAD_425 vpwr_R_branch_5 vpwr_R_425 ${R_R_BUFF}
RP_R_LOAD_426 vpwr_R_branch_6 vpwr_R_426 ${R_R_BUFF}
RP_R_LOAD_427 vpwr_R_branch_0 vpwr_R_427 ${R_R_BUFF}
RP_R_LOAD_428 vpwr_R_branch_1 vpwr_R_428 ${R_R_BUFF}
RP_R_LOAD_429 vpwr_R_branch_2 vpwr_R_429 ${R_R_BUFF}
RP_R_LOAD_430 vpwr_R_branch_3 vpwr_R_430 ${R_R_BUFF}
RP_R_LOAD_431 vpwr_R_branch_4 vpwr_R_431 ${R_R_BUFF}
RP_R_LOAD_432 vpwr_R_branch_5 vpwr_R_432 ${R_R_BUFF}
RP_R_LOAD_433 vpwr_R_branch_6 vpwr_R_433 ${R_R_BUFF}
RP_R_LOAD_434 vpwr_R_branch_0 vpwr_R_434 ${R_R_BUFF}
RP_R_LOAD_435 vpwr_R_branch_1 vpwr_R_435 ${R_R_BUFF}
RP_R_LOAD_436 vpwr_R_branch_2 vpwr_R_436 ${R_R_BUFF}
RP_R_LOAD_437 vpwr_R_branch_3 vpwr_R_437 ${R_R_BUFF}
RP_R_LOAD_438 vpwr_R_branch_4 vpwr_R_438 ${R_R_BUFF}
RP_R_LOAD_439 vpwr_R_branch_5 vpwr_R_439 ${R_R_BUFF}
RP_R_LOAD_440 vpwr_R_branch_6 vpwr_R_440 ${R_R_BUFF}
RP_R_LOAD_441 vpwr_R_branch_0 vpwr_R_441 ${R_R_BUFF}
RP_R_LOAD_442 vpwr_R_branch_1 vpwr_R_442 ${R_R_BUFF}
RP_R_LOAD_443 vpwr_R_branch_2 vpwr_R_443 ${R_R_BUFF}
RP_R_LOAD_444 vpwr_R_branch_3 vpwr_R_444 ${R_R_BUFF}
RP_R_LOAD_445 vpwr_R_branch_4 vpwr_R_445 ${R_R_BUFF}
RP_R_LOAD_446 vpwr_R_branch_5 vpwr_R_446 ${R_R_BUFF}
RP_R_LOAD_447 vpwr_R_branch_6 vpwr_R_447 ${R_R_BUFF}
RP_R_LOAD_448 vpwr_R_branch_0 vpwr_R_448 ${R_R_BUFF}
RP_R_LOAD_449 vpwr_R_branch_1 vpwr_R_449 ${R_R_BUFF}
RP_R_LOAD_450 vpwr_R_branch_2 vpwr_R_450 ${R_R_BUFF}
RP_R_LOAD_451 vpwr_R_branch_3 vpwr_R_451 ${R_R_BUFF}
RP_R_LOAD_452 vpwr_R_branch_4 vpwr_R_452 ${R_R_BUFF}
RP_R_LOAD_453 vpwr_R_branch_5 vpwr_R_453 ${R_R_BUFF}
RP_R_LOAD_454 vpwr_R_branch_6 vpwr_R_454 ${R_R_BUFF}
RP_R_LOAD_455 vpwr_R_branch_0 vpwr_R_455 ${R_R_BUFF}
RP_R_LOAD_456 vpwr_R_branch_1 vpwr_R_456 ${R_R_BUFF}
RP_R_LOAD_457 vpwr_R_branch_2 vpwr_R_457 ${R_R_BUFF}
RP_R_LOAD_458 vpwr_R_branch_3 vpwr_R_458 ${R_R_BUFF}
RP_R_LOAD_459 vpwr_R_branch_4 vpwr_R_459 ${R_R_BUFF}
RP_R_LOAD_460 vpwr_R_branch_5 vpwr_R_460 ${R_R_BUFF}
RP_R_LOAD_461 vpwr_R_branch_6 vpwr_R_461 ${R_R_BUFF}
RP_R_LOAD_462 vpwr_R_branch_0 vpwr_R_462 ${R_R_BUFF}
RP_R_LOAD_463 vpwr_R_branch_1 vpwr_R_463 ${R_R_BUFF}
RP_R_LOAD_464 vpwr_R_branch_2 vpwr_R_464 ${R_R_BUFF}
RP_R_LOAD_465 vpwr_R_branch_3 vpwr_R_465 ${R_R_BUFF}
RP_R_LOAD_466 vpwr_R_branch_4 vpwr_R_466 ${R_R_BUFF}
RP_R_LOAD_467 vpwr_R_branch_5 vpwr_R_467 ${R_R_BUFF}
RP_R_LOAD_468 vpwr_R_branch_6 vpwr_R_468 ${R_R_BUFF}
RP_R_LOAD_469 vpwr_R_branch_0 vpwr_R_469 ${R_R_BUFF}
RP_R_LOAD_470 vpwr_R_branch_1 vpwr_R_470 ${R_R_BUFF}
RP_R_LOAD_471 vpwr_R_branch_2 vpwr_R_471 ${R_R_BUFF}
RP_R_LOAD_472 vpwr_R_branch_3 vpwr_R_472 ${R_R_BUFF}
RP_R_LOAD_473 vpwr_R_branch_4 vpwr_R_473 ${R_R_BUFF}
RP_R_LOAD_474 vpwr_R_branch_5 vpwr_R_474 ${R_R_BUFF}
RP_R_LOAD_475 vpwr_R_branch_6 vpwr_R_475 ${R_R_BUFF}
RP_R_LOAD_476 vpwr_R_branch_0 vpwr_R_476 ${R_R_BUFF}
RP_R_LOAD_477 vpwr_R_branch_1 vpwr_R_477 ${R_R_BUFF}
RP_R_LOAD_478 vpwr_R_branch_2 vpwr_R_478 ${R_R_BUFF}
RP_R_LOAD_479 vpwr_R_branch_3 vpwr_R_479 ${R_R_BUFF}
RP_R_LOAD_480 vpwr_R_branch_4 vpwr_R_480 ${R_R_BUFF}
RP_R_LOAD_481 vpwr_R_branch_5 vpwr_R_481 ${R_R_BUFF}
RP_R_LOAD_482 vpwr_R_branch_6 vpwr_R_482 ${R_R_BUFF}
RP_R_LOAD_483 vpwr_R_branch_0 vpwr_R_483 ${R_R_BUFF}
RP_R_LOAD_484 vpwr_R_branch_1 vpwr_R_484 ${R_R_BUFF}
RP_R_LOAD_485 vpwr_R_branch_2 vpwr_R_485 ${R_R_BUFF}
RP_R_LOAD_486 vpwr_R_branch_3 vpwr_R_486 ${R_R_BUFF}
RP_R_LOAD_487 vpwr_R_branch_4 vpwr_R_487 ${R_R_BUFF}
RP_R_LOAD_488 vpwr_R_branch_5 vpwr_R_488 ${R_R_BUFF}
RP_R_LOAD_489 vpwr_R_branch_6 vpwr_R_489 ${R_R_BUFF}
RP_R_LOAD_490 vpwr_R_branch_0 vpwr_R_490 ${R_R_BUFF}
RP_R_LOAD_491 vpwr_R_branch_1 vpwr_R_491 ${R_R_BUFF}
RP_R_LOAD_492 vpwr_R_branch_2 vpwr_R_492 ${R_R_BUFF}
RP_R_LOAD_493 vpwr_R_branch_3 vpwr_R_493 ${R_R_BUFF}
RP_R_LOAD_494 vpwr_R_branch_4 vpwr_R_494 ${R_R_BUFF}
RP_R_LOAD_495 vpwr_R_branch_5 vpwr_R_495 ${R_R_BUFF}
RP_R_LOAD_496 vpwr_R_branch_6 vpwr_R_496 ${R_R_BUFF}
RP_R_LOAD_497 vpwr_R_branch_0 vpwr_R_497 ${R_R_BUFF}
RP_R_LOAD_498 vpwr_R_branch_1 vpwr_R_498 ${R_R_BUFF}
RP_R_LOAD_499 vpwr_R_branch_2 vpwr_R_499 ${R_R_BUFF}
RP_R_LOAD_500 vpwr_R_branch_3 vpwr_R_500 ${R_R_BUFF}
RP_R_LOAD_501 vpwr_R_branch_4 vpwr_R_501 ${R_R_BUFF}
RP_R_LOAD_502 vpwr_R_branch_5 vpwr_R_502 ${R_R_BUFF}
RP_R_LOAD_503 vpwr_R_branch_6 vpwr_R_503 ${R_R_BUFF}
RP_R_LOAD_504 vpwr_R_branch_0 vpwr_R_504 ${R_R_BUFF}
RP_R_LOAD_505 vpwr_R_branch_1 vpwr_R_505 ${R_R_BUFF}
RP_R_LOAD_506 vpwr_R_branch_2 vpwr_R_506 ${R_R_BUFF}
RP_R_LOAD_507 vpwr_R_branch_3 vpwr_R_507 ${R_R_BUFF}
RP_R_LOAD_508 vpwr_R_branch_4 vpwr_R_508 ${R_R_BUFF}
RP_R_LOAD_509 vpwr_R_branch_5 vpwr_R_509 ${R_R_BUFF}
RP_R_LOAD_510 vpwr_R_branch_6 vpwr_R_510 ${R_R_BUFF}
RP_R_LOAD_511 vpwr_R_branch_0 vpwr_R_511 ${R_R_BUFF}
RP_R_LOAD_512 vpwr_R_branch_1 vpwr_R_512 ${R_R_BUFF}
RP_R_LOAD_513 vpwr_R_branch_2 vpwr_R_513 ${R_R_BUFF}
RP_R_LOAD_514 vpwr_R_branch_3 vpwr_R_514 ${R_R_BUFF}
RP_R_LOAD_515 vpwr_R_branch_4 vpwr_R_515 ${R_R_BUFF}
RP_R_LOAD_516 vpwr_R_branch_5 vpwr_R_516 ${R_R_BUFF}
RP_R_LOAD_517 vpwr_R_branch_6 vpwr_R_517 ${R_R_BUFF}
RP_R_LOAD_518 vpwr_R_branch_0 vpwr_R_518 ${R_R_BUFF}
RP_R_LOAD_519 vpwr_R_branch_1 vpwr_R_519 ${R_R_BUFF}
RP_R_LOAD_520 vpwr_R_branch_2 vpwr_R_520 ${R_R_BUFF}
RP_R_LOAD_521 vpwr_R_branch_3 vpwr_R_521 ${R_R_BUFF}
RP_R_LOAD_522 vpwr_R_branch_4 vpwr_R_522 ${R_R_BUFF}
RP_R_LOAD_523 vpwr_R_branch_5 vpwr_R_523 ${R_R_BUFF}
RP_R_LOAD_524 vpwr_R_branch_6 vpwr_R_524 ${R_R_BUFF}
RP_R_LOAD_525 vpwr_R_branch_0 vpwr_R_525 ${R_R_BUFF}
RP_R_LOAD_526 vpwr_R_branch_1 vpwr_R_526 ${R_R_BUFF}
RP_R_LOAD_527 vpwr_R_branch_2 vpwr_R_527 ${R_R_BUFF}
RP_R_LOAD_528 vpwr_R_branch_3 vpwr_R_528 ${R_R_BUFF}
RP_R_LOAD_529 vpwr_R_branch_4 vpwr_R_529 ${R_R_BUFF}
RP_R_LOAD_530 vpwr_R_branch_5 vpwr_R_530 ${R_R_BUFF}
RP_R_LOAD_531 vpwr_R_branch_6 vpwr_R_531 ${R_R_BUFF}
RP_R_LOAD_532 vpwr_R_branch_0 vpwr_R_532 ${R_R_BUFF}
RP_R_LOAD_533 vpwr_R_branch_1 vpwr_R_533 ${R_R_BUFF}
RP_R_LOAD_534 vpwr_R_branch_2 vpwr_R_534 ${R_R_BUFF}
RP_R_LOAD_535 vpwr_R_branch_3 vpwr_R_535 ${R_R_BUFF}
RP_R_LOAD_536 vpwr_R_branch_4 vpwr_R_536 ${R_R_BUFF}
RP_R_LOAD_537 vpwr_R_branch_5 vpwr_R_537 ${R_R_BUFF}
RP_R_LOAD_538 vpwr_R_branch_6 vpwr_R_538 ${R_R_BUFF}
RP_R_LOAD_539 vpwr_R_branch_0 vpwr_R_539 ${R_R_BUFF}
RP_R_LOAD_540 vpwr_R_branch_1 vpwr_R_540 ${R_R_BUFF}
RP_R_LOAD_541 vpwr_R_branch_2 vpwr_R_541 ${R_R_BUFF}
RP_R_LOAD_542 vpwr_R_branch_3 vpwr_R_542 ${R_R_BUFF}
RP_R_LOAD_543 vpwr_R_branch_4 vpwr_R_543 ${R_R_BUFF}
XDC_R_0_0 VGND VNB vpwr_R_0 vpwr_R_0 sky130_fd_sc_hd__decap_12
XDC_R_1_0 VGND VNB vpwr_R_0 vpwr_R_0 sky130_fd_sc_hd__decap_12
XDC_R_2_0 VGND VNB vpwr_R_0 vpwr_R_0 sky130_fd_sc_hd__decap_12
XDC_R_0_1 VGND VNB vpwr_R_1 vpwr_R_1 sky130_fd_sc_hd__decap_12
XDC_R_1_1 VGND VNB vpwr_R_1 vpwr_R_1 sky130_fd_sc_hd__decap_12
XDC_R_2_1 VGND VNB vpwr_R_1 vpwr_R_1 sky130_fd_sc_hd__decap_12
XDC_R_0_2 VGND VNB vpwr_R_2 vpwr_R_2 sky130_fd_sc_hd__decap_12
XDC_R_1_2 VGND VNB vpwr_R_2 vpwr_R_2 sky130_fd_sc_hd__decap_12
XDC_R_2_2 VGND VNB vpwr_R_2 vpwr_R_2 sky130_fd_sc_hd__decap_12
XDC_R_0_3 VGND VNB vpwr_R_3 vpwr_R_3 sky130_fd_sc_hd__decap_12
XDC_R_1_3 VGND VNB vpwr_R_3 vpwr_R_3 sky130_fd_sc_hd__decap_12
XDC_R_2_3 VGND VNB vpwr_R_3 vpwr_R_3 sky130_fd_sc_hd__decap_12
XDC_R_0_4 VGND VNB vpwr_R_4 vpwr_R_4 sky130_fd_sc_hd__decap_12
XDC_R_1_4 VGND VNB vpwr_R_4 vpwr_R_4 sky130_fd_sc_hd__decap_12
XDC_R_2_4 VGND VNB vpwr_R_4 vpwr_R_4 sky130_fd_sc_hd__decap_12
XDC_R_0_5 VGND VNB vpwr_R_5 vpwr_R_5 sky130_fd_sc_hd__decap_12
XDC_R_1_5 VGND VNB vpwr_R_5 vpwr_R_5 sky130_fd_sc_hd__decap_12
XDC_R_2_5 VGND VNB vpwr_R_5 vpwr_R_5 sky130_fd_sc_hd__decap_12
XDC_R_0_6 VGND VNB vpwr_R_6 vpwr_R_6 sky130_fd_sc_hd__decap_12
XDC_R_1_6 VGND VNB vpwr_R_6 vpwr_R_6 sky130_fd_sc_hd__decap_12
XDC_R_2_6 VGND VNB vpwr_R_6 vpwr_R_6 sky130_fd_sc_hd__decap_12
XDC_R_0_7 VGND VNB vpwr_R_7 vpwr_R_7 sky130_fd_sc_hd__decap_12
XDC_R_1_7 VGND VNB vpwr_R_7 vpwr_R_7 sky130_fd_sc_hd__decap_12
XDC_R_2_7 VGND VNB vpwr_R_7 vpwr_R_7 sky130_fd_sc_hd__decap_12
XDC_R_0_8 VGND VNB vpwr_R_8 vpwr_R_8 sky130_fd_sc_hd__decap_12
XDC_R_1_8 VGND VNB vpwr_R_8 vpwr_R_8 sky130_fd_sc_hd__decap_12
XDC_R_2_8 VGND VNB vpwr_R_8 vpwr_R_8 sky130_fd_sc_hd__decap_12
XDC_R_0_9 VGND VNB vpwr_R_9 vpwr_R_9 sky130_fd_sc_hd__decap_12
XDC_R_1_9 VGND VNB vpwr_R_9 vpwr_R_9 sky130_fd_sc_hd__decap_12
XDC_R_2_9 VGND VNB vpwr_R_9 vpwr_R_9 sky130_fd_sc_hd__decap_12
XDC_R_0_10 VGND VNB vpwr_R_10 vpwr_R_10 sky130_fd_sc_hd__decap_12
XDC_R_1_10 VGND VNB vpwr_R_10 vpwr_R_10 sky130_fd_sc_hd__decap_12
XDC_R_2_10 VGND VNB vpwr_R_10 vpwr_R_10 sky130_fd_sc_hd__decap_12
XDC_R_0_11 VGND VNB vpwr_R_11 vpwr_R_11 sky130_fd_sc_hd__decap_12
XDC_R_1_11 VGND VNB vpwr_R_11 vpwr_R_11 sky130_fd_sc_hd__decap_12
XDC_R_2_11 VGND VNB vpwr_R_11 vpwr_R_11 sky130_fd_sc_hd__decap_12
XDC_R_0_12 VGND VNB vpwr_R_12 vpwr_R_12 sky130_fd_sc_hd__decap_12
XDC_R_1_12 VGND VNB vpwr_R_12 vpwr_R_12 sky130_fd_sc_hd__decap_12
XDC_R_2_12 VGND VNB vpwr_R_12 vpwr_R_12 sky130_fd_sc_hd__decap_12
XDC_R_0_13 VGND VNB vpwr_R_13 vpwr_R_13 sky130_fd_sc_hd__decap_12
XDC_R_1_13 VGND VNB vpwr_R_13 vpwr_R_13 sky130_fd_sc_hd__decap_12
XDC_R_2_13 VGND VNB vpwr_R_13 vpwr_R_13 sky130_fd_sc_hd__decap_12
XDC_R_0_14 VGND VNB vpwr_R_14 vpwr_R_14 sky130_fd_sc_hd__decap_12
XDC_R_1_14 VGND VNB vpwr_R_14 vpwr_R_14 sky130_fd_sc_hd__decap_12
XDC_R_2_14 VGND VNB vpwr_R_14 vpwr_R_14 sky130_fd_sc_hd__decap_12
XDC_R_0_15 VGND VNB vpwr_R_15 vpwr_R_15 sky130_fd_sc_hd__decap_12
XDC_R_1_15 VGND VNB vpwr_R_15 vpwr_R_15 sky130_fd_sc_hd__decap_12
XDC_R_2_15 VGND VNB vpwr_R_15 vpwr_R_15 sky130_fd_sc_hd__decap_12
XDC_R_0_16 VGND VNB vpwr_R_16 vpwr_R_16 sky130_fd_sc_hd__decap_12
XDC_R_1_16 VGND VNB vpwr_R_16 vpwr_R_16 sky130_fd_sc_hd__decap_12
XDC_R_2_16 VGND VNB vpwr_R_16 vpwr_R_16 sky130_fd_sc_hd__decap_12
XDC_R_0_17 VGND VNB vpwr_R_17 vpwr_R_17 sky130_fd_sc_hd__decap_12
XDC_R_1_17 VGND VNB vpwr_R_17 vpwr_R_17 sky130_fd_sc_hd__decap_12
XDC_R_2_17 VGND VNB vpwr_R_17 vpwr_R_17 sky130_fd_sc_hd__decap_12
XDC_R_0_18 VGND VNB vpwr_R_18 vpwr_R_18 sky130_fd_sc_hd__decap_12
XDC_R_1_18 VGND VNB vpwr_R_18 vpwr_R_18 sky130_fd_sc_hd__decap_12
XDC_R_2_18 VGND VNB vpwr_R_18 vpwr_R_18 sky130_fd_sc_hd__decap_12
XDC_R_0_19 VGND VNB vpwr_R_19 vpwr_R_19 sky130_fd_sc_hd__decap_12
XDC_R_1_19 VGND VNB vpwr_R_19 vpwr_R_19 sky130_fd_sc_hd__decap_12
XDC_R_2_19 VGND VNB vpwr_R_19 vpwr_R_19 sky130_fd_sc_hd__decap_12
XDC_R_0_20 VGND VNB vpwr_R_20 vpwr_R_20 sky130_fd_sc_hd__decap_12
XDC_R_1_20 VGND VNB vpwr_R_20 vpwr_R_20 sky130_fd_sc_hd__decap_12
XDC_R_2_20 VGND VNB vpwr_R_20 vpwr_R_20 sky130_fd_sc_hd__decap_12
XDC_R_0_21 VGND VNB vpwr_R_21 vpwr_R_21 sky130_fd_sc_hd__decap_12
XDC_R_1_21 VGND VNB vpwr_R_21 vpwr_R_21 sky130_fd_sc_hd__decap_12
XDC_R_2_21 VGND VNB vpwr_R_21 vpwr_R_21 sky130_fd_sc_hd__decap_12
XDC_R_0_22 VGND VNB vpwr_R_22 vpwr_R_22 sky130_fd_sc_hd__decap_12
XDC_R_1_22 VGND VNB vpwr_R_22 vpwr_R_22 sky130_fd_sc_hd__decap_12
XDC_R_2_22 VGND VNB vpwr_R_22 vpwr_R_22 sky130_fd_sc_hd__decap_12
XDC_R_0_23 VGND VNB vpwr_R_23 vpwr_R_23 sky130_fd_sc_hd__decap_12
XDC_R_1_23 VGND VNB vpwr_R_23 vpwr_R_23 sky130_fd_sc_hd__decap_12
XDC_R_2_23 VGND VNB vpwr_R_23 vpwr_R_23 sky130_fd_sc_hd__decap_12
XDC_R_0_24 VGND VNB vpwr_R_24 vpwr_R_24 sky130_fd_sc_hd__decap_12
XDC_R_1_24 VGND VNB vpwr_R_24 vpwr_R_24 sky130_fd_sc_hd__decap_12
XDC_R_2_24 VGND VNB vpwr_R_24 vpwr_R_24 sky130_fd_sc_hd__decap_12
XDC_R_0_25 VGND VNB vpwr_R_25 vpwr_R_25 sky130_fd_sc_hd__decap_12
XDC_R_1_25 VGND VNB vpwr_R_25 vpwr_R_25 sky130_fd_sc_hd__decap_12
XDC_R_2_25 VGND VNB vpwr_R_25 vpwr_R_25 sky130_fd_sc_hd__decap_12
XDC_R_0_26 VGND VNB vpwr_R_26 vpwr_R_26 sky130_fd_sc_hd__decap_12
XDC_R_1_26 VGND VNB vpwr_R_26 vpwr_R_26 sky130_fd_sc_hd__decap_12
XDC_R_2_26 VGND VNB vpwr_R_26 vpwr_R_26 sky130_fd_sc_hd__decap_12
XDC_R_0_27 VGND VNB vpwr_R_27 vpwr_R_27 sky130_fd_sc_hd__decap_12
XDC_R_1_27 VGND VNB vpwr_R_27 vpwr_R_27 sky130_fd_sc_hd__decap_12
XDC_R_2_27 VGND VNB vpwr_R_27 vpwr_R_27 sky130_fd_sc_hd__decap_12
XDC_R_0_28 VGND VNB vpwr_R_28 vpwr_R_28 sky130_fd_sc_hd__decap_12
XDC_R_1_28 VGND VNB vpwr_R_28 vpwr_R_28 sky130_fd_sc_hd__decap_12
XDC_R_2_28 VGND VNB vpwr_R_28 vpwr_R_28 sky130_fd_sc_hd__decap_12
XDC_R_0_29 VGND VNB vpwr_R_29 vpwr_R_29 sky130_fd_sc_hd__decap_12
XDC_R_1_29 VGND VNB vpwr_R_29 vpwr_R_29 sky130_fd_sc_hd__decap_12
XDC_R_2_29 VGND VNB vpwr_R_29 vpwr_R_29 sky130_fd_sc_hd__decap_12
XDC_R_0_30 VGND VNB vpwr_R_30 vpwr_R_30 sky130_fd_sc_hd__decap_12
XDC_R_1_30 VGND VNB vpwr_R_30 vpwr_R_30 sky130_fd_sc_hd__decap_12
XDC_R_2_30 VGND VNB vpwr_R_30 vpwr_R_30 sky130_fd_sc_hd__decap_12
XDC_R_0_31 VGND VNB vpwr_R_31 vpwr_R_31 sky130_fd_sc_hd__decap_12
XDC_R_1_31 VGND VNB vpwr_R_31 vpwr_R_31 sky130_fd_sc_hd__decap_12
XDC_R_2_31 VGND VNB vpwr_R_31 vpwr_R_31 sky130_fd_sc_hd__decap_12
XDC_R_0_32 VGND VNB vpwr_R_32 vpwr_R_32 sky130_fd_sc_hd__decap_12
XDC_R_1_32 VGND VNB vpwr_R_32 vpwr_R_32 sky130_fd_sc_hd__decap_12
XDC_R_2_32 VGND VNB vpwr_R_32 vpwr_R_32 sky130_fd_sc_hd__decap_12
XDC_R_0_33 VGND VNB vpwr_R_33 vpwr_R_33 sky130_fd_sc_hd__decap_12
XDC_R_1_33 VGND VNB vpwr_R_33 vpwr_R_33 sky130_fd_sc_hd__decap_12
XDC_R_2_33 VGND VNB vpwr_R_33 vpwr_R_33 sky130_fd_sc_hd__decap_12
XDC_R_0_34 VGND VNB vpwr_R_34 vpwr_R_34 sky130_fd_sc_hd__decap_12
XDC_R_1_34 VGND VNB vpwr_R_34 vpwr_R_34 sky130_fd_sc_hd__decap_12
XDC_R_2_34 VGND VNB vpwr_R_34 vpwr_R_34 sky130_fd_sc_hd__decap_12
XDC_R_0_35 VGND VNB vpwr_R_35 vpwr_R_35 sky130_fd_sc_hd__decap_12
XDC_R_1_35 VGND VNB vpwr_R_35 vpwr_R_35 sky130_fd_sc_hd__decap_12
XDC_R_2_35 VGND VNB vpwr_R_35 vpwr_R_35 sky130_fd_sc_hd__decap_12
XDC_R_0_36 VGND VNB vpwr_R_36 vpwr_R_36 sky130_fd_sc_hd__decap_12
XDC_R_1_36 VGND VNB vpwr_R_36 vpwr_R_36 sky130_fd_sc_hd__decap_12
XDC_R_2_36 VGND VNB vpwr_R_36 vpwr_R_36 sky130_fd_sc_hd__decap_12
XDC_R_0_37 VGND VNB vpwr_R_37 vpwr_R_37 sky130_fd_sc_hd__decap_12
XDC_R_1_37 VGND VNB vpwr_R_37 vpwr_R_37 sky130_fd_sc_hd__decap_12
XDC_R_2_37 VGND VNB vpwr_R_37 vpwr_R_37 sky130_fd_sc_hd__decap_12
XDC_R_0_38 VGND VNB vpwr_R_38 vpwr_R_38 sky130_fd_sc_hd__decap_12
XDC_R_1_38 VGND VNB vpwr_R_38 vpwr_R_38 sky130_fd_sc_hd__decap_12
XDC_R_2_38 VGND VNB vpwr_R_38 vpwr_R_38 sky130_fd_sc_hd__decap_12
XDC_R_0_39 VGND VNB vpwr_R_39 vpwr_R_39 sky130_fd_sc_hd__decap_12
XDC_R_1_39 VGND VNB vpwr_R_39 vpwr_R_39 sky130_fd_sc_hd__decap_12
XDC_R_2_39 VGND VNB vpwr_R_39 vpwr_R_39 sky130_fd_sc_hd__decap_12
XDC_R_0_40 VGND VNB vpwr_R_40 vpwr_R_40 sky130_fd_sc_hd__decap_12
XDC_R_1_40 VGND VNB vpwr_R_40 vpwr_R_40 sky130_fd_sc_hd__decap_12
XDC_R_2_40 VGND VNB vpwr_R_40 vpwr_R_40 sky130_fd_sc_hd__decap_12
XDC_R_0_41 VGND VNB vpwr_R_41 vpwr_R_41 sky130_fd_sc_hd__decap_12
XDC_R_1_41 VGND VNB vpwr_R_41 vpwr_R_41 sky130_fd_sc_hd__decap_12
XDC_R_2_41 VGND VNB vpwr_R_41 vpwr_R_41 sky130_fd_sc_hd__decap_12
XDC_R_0_42 VGND VNB vpwr_R_42 vpwr_R_42 sky130_fd_sc_hd__decap_12
XDC_R_1_42 VGND VNB vpwr_R_42 vpwr_R_42 sky130_fd_sc_hd__decap_12
XDC_R_2_42 VGND VNB vpwr_R_42 vpwr_R_42 sky130_fd_sc_hd__decap_12
XDC_R_0_43 VGND VNB vpwr_R_43 vpwr_R_43 sky130_fd_sc_hd__decap_12
XDC_R_1_43 VGND VNB vpwr_R_43 vpwr_R_43 sky130_fd_sc_hd__decap_12
XDC_R_2_43 VGND VNB vpwr_R_43 vpwr_R_43 sky130_fd_sc_hd__decap_12
XDC_R_0_44 VGND VNB vpwr_R_44 vpwr_R_44 sky130_fd_sc_hd__decap_12
XDC_R_1_44 VGND VNB vpwr_R_44 vpwr_R_44 sky130_fd_sc_hd__decap_12
XDC_R_2_44 VGND VNB vpwr_R_44 vpwr_R_44 sky130_fd_sc_hd__decap_12
XDC_R_0_45 VGND VNB vpwr_R_45 vpwr_R_45 sky130_fd_sc_hd__decap_12
XDC_R_1_45 VGND VNB vpwr_R_45 vpwr_R_45 sky130_fd_sc_hd__decap_12
XDC_R_2_45 VGND VNB vpwr_R_45 vpwr_R_45 sky130_fd_sc_hd__decap_12
XDC_R_0_46 VGND VNB vpwr_R_46 vpwr_R_46 sky130_fd_sc_hd__decap_12
XDC_R_1_46 VGND VNB vpwr_R_46 vpwr_R_46 sky130_fd_sc_hd__decap_12
XDC_R_2_46 VGND VNB vpwr_R_46 vpwr_R_46 sky130_fd_sc_hd__decap_12
XDC_R_0_47 VGND VNB vpwr_R_47 vpwr_R_47 sky130_fd_sc_hd__decap_12
XDC_R_1_47 VGND VNB vpwr_R_47 vpwr_R_47 sky130_fd_sc_hd__decap_12
XDC_R_2_47 VGND VNB vpwr_R_47 vpwr_R_47 sky130_fd_sc_hd__decap_12
XDC_R_0_48 VGND VNB vpwr_R_48 vpwr_R_48 sky130_fd_sc_hd__decap_12
XDC_R_1_48 VGND VNB vpwr_R_48 vpwr_R_48 sky130_fd_sc_hd__decap_12
XDC_R_2_48 VGND VNB vpwr_R_48 vpwr_R_48 sky130_fd_sc_hd__decap_12
XDC_R_0_49 VGND VNB vpwr_R_49 vpwr_R_49 sky130_fd_sc_hd__decap_12
XDC_R_1_49 VGND VNB vpwr_R_49 vpwr_R_49 sky130_fd_sc_hd__decap_12
XDC_R_2_49 VGND VNB vpwr_R_49 vpwr_R_49 sky130_fd_sc_hd__decap_12
XDC_R_0_50 VGND VNB vpwr_R_50 vpwr_R_50 sky130_fd_sc_hd__decap_12
XDC_R_1_50 VGND VNB vpwr_R_50 vpwr_R_50 sky130_fd_sc_hd__decap_12
XDC_R_2_50 VGND VNB vpwr_R_50 vpwr_R_50 sky130_fd_sc_hd__decap_12
XDC_R_0_51 VGND VNB vpwr_R_51 vpwr_R_51 sky130_fd_sc_hd__decap_12
XDC_R_1_51 VGND VNB vpwr_R_51 vpwr_R_51 sky130_fd_sc_hd__decap_12
XDC_R_2_51 VGND VNB vpwr_R_51 vpwr_R_51 sky130_fd_sc_hd__decap_12
XDC_R_0_52 VGND VNB vpwr_R_52 vpwr_R_52 sky130_fd_sc_hd__decap_12
XDC_R_1_52 VGND VNB vpwr_R_52 vpwr_R_52 sky130_fd_sc_hd__decap_12
XDC_R_2_52 VGND VNB vpwr_R_52 vpwr_R_52 sky130_fd_sc_hd__decap_12
XDC_R_0_53 VGND VNB vpwr_R_53 vpwr_R_53 sky130_fd_sc_hd__decap_12
XDC_R_1_53 VGND VNB vpwr_R_53 vpwr_R_53 sky130_fd_sc_hd__decap_12
XDC_R_2_53 VGND VNB vpwr_R_53 vpwr_R_53 sky130_fd_sc_hd__decap_12
XDC_R_0_54 VGND VNB vpwr_R_54 vpwr_R_54 sky130_fd_sc_hd__decap_12
XDC_R_1_54 VGND VNB vpwr_R_54 vpwr_R_54 sky130_fd_sc_hd__decap_12
XDC_R_2_54 VGND VNB vpwr_R_54 vpwr_R_54 sky130_fd_sc_hd__decap_12
XDC_R_0_55 VGND VNB vpwr_R_55 vpwr_R_55 sky130_fd_sc_hd__decap_12
XDC_R_1_55 VGND VNB vpwr_R_55 vpwr_R_55 sky130_fd_sc_hd__decap_12
XDC_R_2_55 VGND VNB vpwr_R_55 vpwr_R_55 sky130_fd_sc_hd__decap_12
XDC_R_0_56 VGND VNB vpwr_R_56 vpwr_R_56 sky130_fd_sc_hd__decap_12
XDC_R_1_56 VGND VNB vpwr_R_56 vpwr_R_56 sky130_fd_sc_hd__decap_12
XDC_R_2_56 VGND VNB vpwr_R_56 vpwr_R_56 sky130_fd_sc_hd__decap_12
XDC_R_0_57 VGND VNB vpwr_R_57 vpwr_R_57 sky130_fd_sc_hd__decap_12
XDC_R_1_57 VGND VNB vpwr_R_57 vpwr_R_57 sky130_fd_sc_hd__decap_12
XDC_R_2_57 VGND VNB vpwr_R_57 vpwr_R_57 sky130_fd_sc_hd__decap_12
XDC_R_0_58 VGND VNB vpwr_R_58 vpwr_R_58 sky130_fd_sc_hd__decap_12
XDC_R_1_58 VGND VNB vpwr_R_58 vpwr_R_58 sky130_fd_sc_hd__decap_12
XDC_R_2_58 VGND VNB vpwr_R_58 vpwr_R_58 sky130_fd_sc_hd__decap_12
XDC_R_0_59 VGND VNB vpwr_R_59 vpwr_R_59 sky130_fd_sc_hd__decap_12
XDC_R_1_59 VGND VNB vpwr_R_59 vpwr_R_59 sky130_fd_sc_hd__decap_12
XDC_R_2_59 VGND VNB vpwr_R_59 vpwr_R_59 sky130_fd_sc_hd__decap_12
XDC_R_0_60 VGND VNB vpwr_R_60 vpwr_R_60 sky130_fd_sc_hd__decap_12
XDC_R_1_60 VGND VNB vpwr_R_60 vpwr_R_60 sky130_fd_sc_hd__decap_12
XDC_R_2_60 VGND VNB vpwr_R_60 vpwr_R_60 sky130_fd_sc_hd__decap_12
XDC_R_0_61 VGND VNB vpwr_R_61 vpwr_R_61 sky130_fd_sc_hd__decap_12
XDC_R_1_61 VGND VNB vpwr_R_61 vpwr_R_61 sky130_fd_sc_hd__decap_12
XDC_R_2_61 VGND VNB vpwr_R_61 vpwr_R_61 sky130_fd_sc_hd__decap_12
XDC_R_0_62 VGND VNB vpwr_R_62 vpwr_R_62 sky130_fd_sc_hd__decap_12
XDC_R_1_62 VGND VNB vpwr_R_62 vpwr_R_62 sky130_fd_sc_hd__decap_12
XDC_R_2_62 VGND VNB vpwr_R_62 vpwr_R_62 sky130_fd_sc_hd__decap_12
XDC_R_0_63 VGND VNB vpwr_R_63 vpwr_R_63 sky130_fd_sc_hd__decap_12
XDC_R_1_63 VGND VNB vpwr_R_63 vpwr_R_63 sky130_fd_sc_hd__decap_12
XDC_R_2_63 VGND VNB vpwr_R_63 vpwr_R_63 sky130_fd_sc_hd__decap_12
XDC_R_0_64 VGND VNB vpwr_R_64 vpwr_R_64 sky130_fd_sc_hd__decap_12
XDC_R_1_64 VGND VNB vpwr_R_64 vpwr_R_64 sky130_fd_sc_hd__decap_12
XDC_R_2_64 VGND VNB vpwr_R_64 vpwr_R_64 sky130_fd_sc_hd__decap_12
XDC_R_0_65 VGND VNB vpwr_R_65 vpwr_R_65 sky130_fd_sc_hd__decap_12
XDC_R_1_65 VGND VNB vpwr_R_65 vpwr_R_65 sky130_fd_sc_hd__decap_12
XDC_R_2_65 VGND VNB vpwr_R_65 vpwr_R_65 sky130_fd_sc_hd__decap_12
XDC_R_0_66 VGND VNB vpwr_R_66 vpwr_R_66 sky130_fd_sc_hd__decap_12
XDC_R_1_66 VGND VNB vpwr_R_66 vpwr_R_66 sky130_fd_sc_hd__decap_12
XDC_R_2_66 VGND VNB vpwr_R_66 vpwr_R_66 sky130_fd_sc_hd__decap_12
XDC_R_0_67 VGND VNB vpwr_R_67 vpwr_R_67 sky130_fd_sc_hd__decap_12
XDC_R_1_67 VGND VNB vpwr_R_67 vpwr_R_67 sky130_fd_sc_hd__decap_12
XDC_R_2_67 VGND VNB vpwr_R_67 vpwr_R_67 sky130_fd_sc_hd__decap_12
XDC_R_0_68 VGND VNB vpwr_R_68 vpwr_R_68 sky130_fd_sc_hd__decap_12
XDC_R_1_68 VGND VNB vpwr_R_68 vpwr_R_68 sky130_fd_sc_hd__decap_12
XDC_R_2_68 VGND VNB vpwr_R_68 vpwr_R_68 sky130_fd_sc_hd__decap_12
XDC_R_0_69 VGND VNB vpwr_R_69 vpwr_R_69 sky130_fd_sc_hd__decap_12
XDC_R_1_69 VGND VNB vpwr_R_69 vpwr_R_69 sky130_fd_sc_hd__decap_12
XDC_R_2_69 VGND VNB vpwr_R_69 vpwr_R_69 sky130_fd_sc_hd__decap_12
XDC_R_0_70 VGND VNB vpwr_R_70 vpwr_R_70 sky130_fd_sc_hd__decap_12
XDC_R_1_70 VGND VNB vpwr_R_70 vpwr_R_70 sky130_fd_sc_hd__decap_12
XDC_R_2_70 VGND VNB vpwr_R_70 vpwr_R_70 sky130_fd_sc_hd__decap_12
XDC_R_0_71 VGND VNB vpwr_R_71 vpwr_R_71 sky130_fd_sc_hd__decap_12
XDC_R_1_71 VGND VNB vpwr_R_71 vpwr_R_71 sky130_fd_sc_hd__decap_12
XDC_R_2_71 VGND VNB vpwr_R_71 vpwr_R_71 sky130_fd_sc_hd__decap_12
XDC_R_0_72 VGND VNB vpwr_R_72 vpwr_R_72 sky130_fd_sc_hd__decap_12
XDC_R_1_72 VGND VNB vpwr_R_72 vpwr_R_72 sky130_fd_sc_hd__decap_12
XDC_R_2_72 VGND VNB vpwr_R_72 vpwr_R_72 sky130_fd_sc_hd__decap_12
XDC_R_0_73 VGND VNB vpwr_R_73 vpwr_R_73 sky130_fd_sc_hd__decap_12
XDC_R_1_73 VGND VNB vpwr_R_73 vpwr_R_73 sky130_fd_sc_hd__decap_12
XDC_R_2_73 VGND VNB vpwr_R_73 vpwr_R_73 sky130_fd_sc_hd__decap_12
XDC_R_0_74 VGND VNB vpwr_R_74 vpwr_R_74 sky130_fd_sc_hd__decap_12
XDC_R_1_74 VGND VNB vpwr_R_74 vpwr_R_74 sky130_fd_sc_hd__decap_12
XDC_R_2_74 VGND VNB vpwr_R_74 vpwr_R_74 sky130_fd_sc_hd__decap_12
XDC_R_0_75 VGND VNB vpwr_R_75 vpwr_R_75 sky130_fd_sc_hd__decap_12
XDC_R_1_75 VGND VNB vpwr_R_75 vpwr_R_75 sky130_fd_sc_hd__decap_12
XDC_R_2_75 VGND VNB vpwr_R_75 vpwr_R_75 sky130_fd_sc_hd__decap_12
XDC_R_0_76 VGND VNB vpwr_R_76 vpwr_R_76 sky130_fd_sc_hd__decap_12
XDC_R_1_76 VGND VNB vpwr_R_76 vpwr_R_76 sky130_fd_sc_hd__decap_12
XDC_R_2_76 VGND VNB vpwr_R_76 vpwr_R_76 sky130_fd_sc_hd__decap_12
XDC_R_0_77 VGND VNB vpwr_R_77 vpwr_R_77 sky130_fd_sc_hd__decap_12
XDC_R_1_77 VGND VNB vpwr_R_77 vpwr_R_77 sky130_fd_sc_hd__decap_12
XDC_R_2_77 VGND VNB vpwr_R_77 vpwr_R_77 sky130_fd_sc_hd__decap_12
XDC_R_0_78 VGND VNB vpwr_R_78 vpwr_R_78 sky130_fd_sc_hd__decap_12
XDC_R_1_78 VGND VNB vpwr_R_78 vpwr_R_78 sky130_fd_sc_hd__decap_12
XDC_R_2_78 VGND VNB vpwr_R_78 vpwr_R_78 sky130_fd_sc_hd__decap_12
XDC_R_0_79 VGND VNB vpwr_R_79 vpwr_R_79 sky130_fd_sc_hd__decap_12
XDC_R_1_79 VGND VNB vpwr_R_79 vpwr_R_79 sky130_fd_sc_hd__decap_12
XDC_R_2_79 VGND VNB vpwr_R_79 vpwr_R_79 sky130_fd_sc_hd__decap_12
XDC_R_0_80 VGND VNB vpwr_R_80 vpwr_R_80 sky130_fd_sc_hd__decap_12
XDC_R_1_80 VGND VNB vpwr_R_80 vpwr_R_80 sky130_fd_sc_hd__decap_12
XDC_R_2_80 VGND VNB vpwr_R_80 vpwr_R_80 sky130_fd_sc_hd__decap_12
XDC_R_0_81 VGND VNB vpwr_R_81 vpwr_R_81 sky130_fd_sc_hd__decap_12
XDC_R_1_81 VGND VNB vpwr_R_81 vpwr_R_81 sky130_fd_sc_hd__decap_12
XDC_R_2_81 VGND VNB vpwr_R_81 vpwr_R_81 sky130_fd_sc_hd__decap_12
XDC_R_0_82 VGND VNB vpwr_R_82 vpwr_R_82 sky130_fd_sc_hd__decap_12
XDC_R_1_82 VGND VNB vpwr_R_82 vpwr_R_82 sky130_fd_sc_hd__decap_12
XDC_R_2_82 VGND VNB vpwr_R_82 vpwr_R_82 sky130_fd_sc_hd__decap_12
XDC_R_0_83 VGND VNB vpwr_R_83 vpwr_R_83 sky130_fd_sc_hd__decap_12
XDC_R_1_83 VGND VNB vpwr_R_83 vpwr_R_83 sky130_fd_sc_hd__decap_12
XDC_R_2_83 VGND VNB vpwr_R_83 vpwr_R_83 sky130_fd_sc_hd__decap_12
XDC_R_0_84 VGND VNB vpwr_R_84 vpwr_R_84 sky130_fd_sc_hd__decap_12
XDC_R_1_84 VGND VNB vpwr_R_84 vpwr_R_84 sky130_fd_sc_hd__decap_12
XDC_R_2_84 VGND VNB vpwr_R_84 vpwr_R_84 sky130_fd_sc_hd__decap_12
XDC_R_0_85 VGND VNB vpwr_R_85 vpwr_R_85 sky130_fd_sc_hd__decap_12
XDC_R_1_85 VGND VNB vpwr_R_85 vpwr_R_85 sky130_fd_sc_hd__decap_12
XDC_R_2_85 VGND VNB vpwr_R_85 vpwr_R_85 sky130_fd_sc_hd__decap_12
XDC_R_0_86 VGND VNB vpwr_R_86 vpwr_R_86 sky130_fd_sc_hd__decap_12
XDC_R_1_86 VGND VNB vpwr_R_86 vpwr_R_86 sky130_fd_sc_hd__decap_12
XDC_R_2_86 VGND VNB vpwr_R_86 vpwr_R_86 sky130_fd_sc_hd__decap_12
XDC_R_0_87 VGND VNB vpwr_R_87 vpwr_R_87 sky130_fd_sc_hd__decap_12
XDC_R_1_87 VGND VNB vpwr_R_87 vpwr_R_87 sky130_fd_sc_hd__decap_12
XDC_R_2_87 VGND VNB vpwr_R_87 vpwr_R_87 sky130_fd_sc_hd__decap_12
XDC_R_0_88 VGND VNB vpwr_R_88 vpwr_R_88 sky130_fd_sc_hd__decap_12
XDC_R_1_88 VGND VNB vpwr_R_88 vpwr_R_88 sky130_fd_sc_hd__decap_12
XDC_R_2_88 VGND VNB vpwr_R_88 vpwr_R_88 sky130_fd_sc_hd__decap_12
XDC_R_0_89 VGND VNB vpwr_R_89 vpwr_R_89 sky130_fd_sc_hd__decap_12
XDC_R_1_89 VGND VNB vpwr_R_89 vpwr_R_89 sky130_fd_sc_hd__decap_12
XDC_R_2_89 VGND VNB vpwr_R_89 vpwr_R_89 sky130_fd_sc_hd__decap_12
XDC_R_0_90 VGND VNB vpwr_R_90 vpwr_R_90 sky130_fd_sc_hd__decap_12
XDC_R_1_90 VGND VNB vpwr_R_90 vpwr_R_90 sky130_fd_sc_hd__decap_12
XDC_R_2_90 VGND VNB vpwr_R_90 vpwr_R_90 sky130_fd_sc_hd__decap_12
XDC_R_0_91 VGND VNB vpwr_R_91 vpwr_R_91 sky130_fd_sc_hd__decap_12
XDC_R_1_91 VGND VNB vpwr_R_91 vpwr_R_91 sky130_fd_sc_hd__decap_12
XDC_R_2_91 VGND VNB vpwr_R_91 vpwr_R_91 sky130_fd_sc_hd__decap_12
XDC_R_0_92 VGND VNB vpwr_R_92 vpwr_R_92 sky130_fd_sc_hd__decap_12
XDC_R_1_92 VGND VNB vpwr_R_92 vpwr_R_92 sky130_fd_sc_hd__decap_12
XDC_R_2_92 VGND VNB vpwr_R_92 vpwr_R_92 sky130_fd_sc_hd__decap_12
XDC_R_0_93 VGND VNB vpwr_R_93 vpwr_R_93 sky130_fd_sc_hd__decap_12
XDC_R_1_93 VGND VNB vpwr_R_93 vpwr_R_93 sky130_fd_sc_hd__decap_12
XDC_R_2_93 VGND VNB vpwr_R_93 vpwr_R_93 sky130_fd_sc_hd__decap_12
XDC_R_0_94 VGND VNB vpwr_R_94 vpwr_R_94 sky130_fd_sc_hd__decap_12
XDC_R_1_94 VGND VNB vpwr_R_94 vpwr_R_94 sky130_fd_sc_hd__decap_12
XDC_R_2_94 VGND VNB vpwr_R_94 vpwr_R_94 sky130_fd_sc_hd__decap_12
XDC_R_0_95 VGND VNB vpwr_R_95 vpwr_R_95 sky130_fd_sc_hd__decap_12
XDC_R_1_95 VGND VNB vpwr_R_95 vpwr_R_95 sky130_fd_sc_hd__decap_12
XDC_R_2_95 VGND VNB vpwr_R_95 vpwr_R_95 sky130_fd_sc_hd__decap_12
XDC_R_0_96 VGND VNB vpwr_R_96 vpwr_R_96 sky130_fd_sc_hd__decap_12
XDC_R_1_96 VGND VNB vpwr_R_96 vpwr_R_96 sky130_fd_sc_hd__decap_12
XDC_R_2_96 VGND VNB vpwr_R_96 vpwr_R_96 sky130_fd_sc_hd__decap_12
XDC_R_0_97 VGND VNB vpwr_R_97 vpwr_R_97 sky130_fd_sc_hd__decap_12
XDC_R_1_97 VGND VNB vpwr_R_97 vpwr_R_97 sky130_fd_sc_hd__decap_12
XDC_R_2_97 VGND VNB vpwr_R_97 vpwr_R_97 sky130_fd_sc_hd__decap_12
XDC_R_0_98 VGND VNB vpwr_R_98 vpwr_R_98 sky130_fd_sc_hd__decap_12
XDC_R_1_98 VGND VNB vpwr_R_98 vpwr_R_98 sky130_fd_sc_hd__decap_12
XDC_R_2_98 VGND VNB vpwr_R_98 vpwr_R_98 sky130_fd_sc_hd__decap_12
XDC_R_0_99 VGND VNB vpwr_R_99 vpwr_R_99 sky130_fd_sc_hd__decap_12
XDC_R_1_99 VGND VNB vpwr_R_99 vpwr_R_99 sky130_fd_sc_hd__decap_12
XDC_R_2_99 VGND VNB vpwr_R_99 vpwr_R_99 sky130_fd_sc_hd__decap_12
XDC_R_0_100 VGND VNB vpwr_R_100 vpwr_R_100 sky130_fd_sc_hd__decap_12
XDC_R_1_100 VGND VNB vpwr_R_100 vpwr_R_100 sky130_fd_sc_hd__decap_12
XDC_R_2_100 VGND VNB vpwr_R_100 vpwr_R_100 sky130_fd_sc_hd__decap_12
XDC_R_0_101 VGND VNB vpwr_R_101 vpwr_R_101 sky130_fd_sc_hd__decap_12
XDC_R_1_101 VGND VNB vpwr_R_101 vpwr_R_101 sky130_fd_sc_hd__decap_12
XDC_R_2_101 VGND VNB vpwr_R_101 vpwr_R_101 sky130_fd_sc_hd__decap_12
XDC_R_0_102 VGND VNB vpwr_R_102 vpwr_R_102 sky130_fd_sc_hd__decap_12
XDC_R_1_102 VGND VNB vpwr_R_102 vpwr_R_102 sky130_fd_sc_hd__decap_12
XDC_R_2_102 VGND VNB vpwr_R_102 vpwr_R_102 sky130_fd_sc_hd__decap_12
XDC_R_0_103 VGND VNB vpwr_R_103 vpwr_R_103 sky130_fd_sc_hd__decap_12
XDC_R_1_103 VGND VNB vpwr_R_103 vpwr_R_103 sky130_fd_sc_hd__decap_12
XDC_R_2_103 VGND VNB vpwr_R_103 vpwr_R_103 sky130_fd_sc_hd__decap_12
XDC_R_0_104 VGND VNB vpwr_R_104 vpwr_R_104 sky130_fd_sc_hd__decap_12
XDC_R_1_104 VGND VNB vpwr_R_104 vpwr_R_104 sky130_fd_sc_hd__decap_12
XDC_R_2_104 VGND VNB vpwr_R_104 vpwr_R_104 sky130_fd_sc_hd__decap_12
XDC_R_0_105 VGND VNB vpwr_R_105 vpwr_R_105 sky130_fd_sc_hd__decap_12
XDC_R_1_105 VGND VNB vpwr_R_105 vpwr_R_105 sky130_fd_sc_hd__decap_12
XDC_R_2_105 VGND VNB vpwr_R_105 vpwr_R_105 sky130_fd_sc_hd__decap_12
XDC_R_0_106 VGND VNB vpwr_R_106 vpwr_R_106 sky130_fd_sc_hd__decap_12
XDC_R_1_106 VGND VNB vpwr_R_106 vpwr_R_106 sky130_fd_sc_hd__decap_12
XDC_R_2_106 VGND VNB vpwr_R_106 vpwr_R_106 sky130_fd_sc_hd__decap_12
XDC_R_0_107 VGND VNB vpwr_R_107 vpwr_R_107 sky130_fd_sc_hd__decap_12
XDC_R_1_107 VGND VNB vpwr_R_107 vpwr_R_107 sky130_fd_sc_hd__decap_12
XDC_R_2_107 VGND VNB vpwr_R_107 vpwr_R_107 sky130_fd_sc_hd__decap_12
XDC_R_0_108 VGND VNB vpwr_R_108 vpwr_R_108 sky130_fd_sc_hd__decap_12
XDC_R_1_108 VGND VNB vpwr_R_108 vpwr_R_108 sky130_fd_sc_hd__decap_12
XDC_R_2_108 VGND VNB vpwr_R_108 vpwr_R_108 sky130_fd_sc_hd__decap_12
XDC_R_0_109 VGND VNB vpwr_R_109 vpwr_R_109 sky130_fd_sc_hd__decap_12
XDC_R_1_109 VGND VNB vpwr_R_109 vpwr_R_109 sky130_fd_sc_hd__decap_12
XDC_R_2_109 VGND VNB vpwr_R_109 vpwr_R_109 sky130_fd_sc_hd__decap_12
XDC_R_0_110 VGND VNB vpwr_R_110 vpwr_R_110 sky130_fd_sc_hd__decap_12
XDC_R_1_110 VGND VNB vpwr_R_110 vpwr_R_110 sky130_fd_sc_hd__decap_12
XDC_R_2_110 VGND VNB vpwr_R_110 vpwr_R_110 sky130_fd_sc_hd__decap_12
XDC_R_0_111 VGND VNB vpwr_R_111 vpwr_R_111 sky130_fd_sc_hd__decap_12
XDC_R_1_111 VGND VNB vpwr_R_111 vpwr_R_111 sky130_fd_sc_hd__decap_12
XDC_R_2_111 VGND VNB vpwr_R_111 vpwr_R_111 sky130_fd_sc_hd__decap_12
XDC_R_0_112 VGND VNB vpwr_R_112 vpwr_R_112 sky130_fd_sc_hd__decap_12
XDC_R_1_112 VGND VNB vpwr_R_112 vpwr_R_112 sky130_fd_sc_hd__decap_12
XDC_R_2_112 VGND VNB vpwr_R_112 vpwr_R_112 sky130_fd_sc_hd__decap_12
XDC_R_0_113 VGND VNB vpwr_R_113 vpwr_R_113 sky130_fd_sc_hd__decap_12
XDC_R_1_113 VGND VNB vpwr_R_113 vpwr_R_113 sky130_fd_sc_hd__decap_12
XDC_R_2_113 VGND VNB vpwr_R_113 vpwr_R_113 sky130_fd_sc_hd__decap_12
XDC_R_0_114 VGND VNB vpwr_R_114 vpwr_R_114 sky130_fd_sc_hd__decap_12
XDC_R_1_114 VGND VNB vpwr_R_114 vpwr_R_114 sky130_fd_sc_hd__decap_12
XDC_R_2_114 VGND VNB vpwr_R_114 vpwr_R_114 sky130_fd_sc_hd__decap_12
XDC_R_0_115 VGND VNB vpwr_R_115 vpwr_R_115 sky130_fd_sc_hd__decap_12
XDC_R_1_115 VGND VNB vpwr_R_115 vpwr_R_115 sky130_fd_sc_hd__decap_12
XDC_R_2_115 VGND VNB vpwr_R_115 vpwr_R_115 sky130_fd_sc_hd__decap_12
XDC_R_0_116 VGND VNB vpwr_R_116 vpwr_R_116 sky130_fd_sc_hd__decap_12
XDC_R_1_116 VGND VNB vpwr_R_116 vpwr_R_116 sky130_fd_sc_hd__decap_12
XDC_R_2_116 VGND VNB vpwr_R_116 vpwr_R_116 sky130_fd_sc_hd__decap_12
XDC_R_0_117 VGND VNB vpwr_R_117 vpwr_R_117 sky130_fd_sc_hd__decap_12
XDC_R_1_117 VGND VNB vpwr_R_117 vpwr_R_117 sky130_fd_sc_hd__decap_12
XDC_R_2_117 VGND VNB vpwr_R_117 vpwr_R_117 sky130_fd_sc_hd__decap_12
XDC_R_0_118 VGND VNB vpwr_R_118 vpwr_R_118 sky130_fd_sc_hd__decap_12
XDC_R_1_118 VGND VNB vpwr_R_118 vpwr_R_118 sky130_fd_sc_hd__decap_12
XDC_R_2_118 VGND VNB vpwr_R_118 vpwr_R_118 sky130_fd_sc_hd__decap_12
XDC_R_0_119 VGND VNB vpwr_R_119 vpwr_R_119 sky130_fd_sc_hd__decap_12
XDC_R_1_119 VGND VNB vpwr_R_119 vpwr_R_119 sky130_fd_sc_hd__decap_12
XDC_R_2_119 VGND VNB vpwr_R_119 vpwr_R_119 sky130_fd_sc_hd__decap_12
XDC_R_0_120 VGND VNB vpwr_R_120 vpwr_R_120 sky130_fd_sc_hd__decap_12
XDC_R_1_120 VGND VNB vpwr_R_120 vpwr_R_120 sky130_fd_sc_hd__decap_12
XDC_R_2_120 VGND VNB vpwr_R_120 vpwr_R_120 sky130_fd_sc_hd__decap_12
XDC_R_0_121 VGND VNB vpwr_R_121 vpwr_R_121 sky130_fd_sc_hd__decap_12
XDC_R_1_121 VGND VNB vpwr_R_121 vpwr_R_121 sky130_fd_sc_hd__decap_12
XDC_R_2_121 VGND VNB vpwr_R_121 vpwr_R_121 sky130_fd_sc_hd__decap_12
XDC_R_0_122 VGND VNB vpwr_R_122 vpwr_R_122 sky130_fd_sc_hd__decap_12
XDC_R_1_122 VGND VNB vpwr_R_122 vpwr_R_122 sky130_fd_sc_hd__decap_12
XDC_R_2_122 VGND VNB vpwr_R_122 vpwr_R_122 sky130_fd_sc_hd__decap_12
XDC_R_0_123 VGND VNB vpwr_R_123 vpwr_R_123 sky130_fd_sc_hd__decap_12
XDC_R_1_123 VGND VNB vpwr_R_123 vpwr_R_123 sky130_fd_sc_hd__decap_12
XDC_R_2_123 VGND VNB vpwr_R_123 vpwr_R_123 sky130_fd_sc_hd__decap_12
XDC_R_0_124 VGND VNB vpwr_R_124 vpwr_R_124 sky130_fd_sc_hd__decap_12
XDC_R_1_124 VGND VNB vpwr_R_124 vpwr_R_124 sky130_fd_sc_hd__decap_12
XDC_R_2_124 VGND VNB vpwr_R_124 vpwr_R_124 sky130_fd_sc_hd__decap_12
XDC_R_0_125 VGND VNB vpwr_R_125 vpwr_R_125 sky130_fd_sc_hd__decap_12
XDC_R_1_125 VGND VNB vpwr_R_125 vpwr_R_125 sky130_fd_sc_hd__decap_12
XDC_R_2_125 VGND VNB vpwr_R_125 vpwr_R_125 sky130_fd_sc_hd__decap_12
XDC_R_0_126 VGND VNB vpwr_R_126 vpwr_R_126 sky130_fd_sc_hd__decap_12
XDC_R_1_126 VGND VNB vpwr_R_126 vpwr_R_126 sky130_fd_sc_hd__decap_12
XDC_R_2_126 VGND VNB vpwr_R_126 vpwr_R_126 sky130_fd_sc_hd__decap_12
XDC_R_0_127 VGND VNB vpwr_R_127 vpwr_R_127 sky130_fd_sc_hd__decap_12
XDC_R_1_127 VGND VNB vpwr_R_127 vpwr_R_127 sky130_fd_sc_hd__decap_12
XDC_R_2_127 VGND VNB vpwr_R_127 vpwr_R_127 sky130_fd_sc_hd__decap_12
XDC_R_0_128 VGND VNB vpwr_R_128 vpwr_R_128 sky130_fd_sc_hd__decap_12
XDC_R_1_128 VGND VNB vpwr_R_128 vpwr_R_128 sky130_fd_sc_hd__decap_12
XDC_R_2_128 VGND VNB vpwr_R_128 vpwr_R_128 sky130_fd_sc_hd__decap_12
XDC_R_0_129 VGND VNB vpwr_R_129 vpwr_R_129 sky130_fd_sc_hd__decap_12
XDC_R_1_129 VGND VNB vpwr_R_129 vpwr_R_129 sky130_fd_sc_hd__decap_12
XDC_R_2_129 VGND VNB vpwr_R_129 vpwr_R_129 sky130_fd_sc_hd__decap_12
XDC_R_0_130 VGND VNB vpwr_R_130 vpwr_R_130 sky130_fd_sc_hd__decap_12
XDC_R_1_130 VGND VNB vpwr_R_130 vpwr_R_130 sky130_fd_sc_hd__decap_12
XDC_R_2_130 VGND VNB vpwr_R_130 vpwr_R_130 sky130_fd_sc_hd__decap_12
XDC_R_0_131 VGND VNB vpwr_R_131 vpwr_R_131 sky130_fd_sc_hd__decap_12
XDC_R_1_131 VGND VNB vpwr_R_131 vpwr_R_131 sky130_fd_sc_hd__decap_12
XDC_R_2_131 VGND VNB vpwr_R_131 vpwr_R_131 sky130_fd_sc_hd__decap_12
XDC_R_0_132 VGND VNB vpwr_R_132 vpwr_R_132 sky130_fd_sc_hd__decap_12
XDC_R_1_132 VGND VNB vpwr_R_132 vpwr_R_132 sky130_fd_sc_hd__decap_12
XDC_R_2_132 VGND VNB vpwr_R_132 vpwr_R_132 sky130_fd_sc_hd__decap_12
XDC_R_0_133 VGND VNB vpwr_R_133 vpwr_R_133 sky130_fd_sc_hd__decap_12
XDC_R_1_133 VGND VNB vpwr_R_133 vpwr_R_133 sky130_fd_sc_hd__decap_12
XDC_R_2_133 VGND VNB vpwr_R_133 vpwr_R_133 sky130_fd_sc_hd__decap_12
XDC_R_0_134 VGND VNB vpwr_R_134 vpwr_R_134 sky130_fd_sc_hd__decap_12
XDC_R_1_134 VGND VNB vpwr_R_134 vpwr_R_134 sky130_fd_sc_hd__decap_12
XDC_R_2_134 VGND VNB vpwr_R_134 vpwr_R_134 sky130_fd_sc_hd__decap_12
XDC_R_0_135 VGND VNB vpwr_R_135 vpwr_R_135 sky130_fd_sc_hd__decap_12
XDC_R_1_135 VGND VNB vpwr_R_135 vpwr_R_135 sky130_fd_sc_hd__decap_12
XDC_R_2_135 VGND VNB vpwr_R_135 vpwr_R_135 sky130_fd_sc_hd__decap_12
XDC_R_0_136 VGND VNB vpwr_R_136 vpwr_R_136 sky130_fd_sc_hd__decap_12
XDC_R_1_136 VGND VNB vpwr_R_136 vpwr_R_136 sky130_fd_sc_hd__decap_12
XDC_R_2_136 VGND VNB vpwr_R_136 vpwr_R_136 sky130_fd_sc_hd__decap_12
XDC_R_0_137 VGND VNB vpwr_R_137 vpwr_R_137 sky130_fd_sc_hd__decap_12
XDC_R_1_137 VGND VNB vpwr_R_137 vpwr_R_137 sky130_fd_sc_hd__decap_12
XDC_R_2_137 VGND VNB vpwr_R_137 vpwr_R_137 sky130_fd_sc_hd__decap_12
XDC_R_0_138 VGND VNB vpwr_R_138 vpwr_R_138 sky130_fd_sc_hd__decap_12
XDC_R_1_138 VGND VNB vpwr_R_138 vpwr_R_138 sky130_fd_sc_hd__decap_12
XDC_R_2_138 VGND VNB vpwr_R_138 vpwr_R_138 sky130_fd_sc_hd__decap_12
XDC_R_0_139 VGND VNB vpwr_R_139 vpwr_R_139 sky130_fd_sc_hd__decap_12
XDC_R_1_139 VGND VNB vpwr_R_139 vpwr_R_139 sky130_fd_sc_hd__decap_12
XDC_R_2_139 VGND VNB vpwr_R_139 vpwr_R_139 sky130_fd_sc_hd__decap_12
XDC_R_0_140 VGND VNB vpwr_R_140 vpwr_R_140 sky130_fd_sc_hd__decap_12
XDC_R_1_140 VGND VNB vpwr_R_140 vpwr_R_140 sky130_fd_sc_hd__decap_12
XDC_R_2_140 VGND VNB vpwr_R_140 vpwr_R_140 sky130_fd_sc_hd__decap_12
XDC_R_0_141 VGND VNB vpwr_R_141 vpwr_R_141 sky130_fd_sc_hd__decap_12
XDC_R_1_141 VGND VNB vpwr_R_141 vpwr_R_141 sky130_fd_sc_hd__decap_12
XDC_R_2_141 VGND VNB vpwr_R_141 vpwr_R_141 sky130_fd_sc_hd__decap_12
XDC_R_0_142 VGND VNB vpwr_R_142 vpwr_R_142 sky130_fd_sc_hd__decap_12
XDC_R_1_142 VGND VNB vpwr_R_142 vpwr_R_142 sky130_fd_sc_hd__decap_12
XDC_R_2_142 VGND VNB vpwr_R_142 vpwr_R_142 sky130_fd_sc_hd__decap_12
XDC_R_0_143 VGND VNB vpwr_R_143 vpwr_R_143 sky130_fd_sc_hd__decap_12
XDC_R_1_143 VGND VNB vpwr_R_143 vpwr_R_143 sky130_fd_sc_hd__decap_12
XDC_R_2_143 VGND VNB vpwr_R_143 vpwr_R_143 sky130_fd_sc_hd__decap_12
XDC_R_0_144 VGND VNB vpwr_R_144 vpwr_R_144 sky130_fd_sc_hd__decap_12
XDC_R_1_144 VGND VNB vpwr_R_144 vpwr_R_144 sky130_fd_sc_hd__decap_12
XDC_R_2_144 VGND VNB vpwr_R_144 vpwr_R_144 sky130_fd_sc_hd__decap_12
XDC_R_0_145 VGND VNB vpwr_R_145 vpwr_R_145 sky130_fd_sc_hd__decap_12
XDC_R_1_145 VGND VNB vpwr_R_145 vpwr_R_145 sky130_fd_sc_hd__decap_12
XDC_R_2_145 VGND VNB vpwr_R_145 vpwr_R_145 sky130_fd_sc_hd__decap_12
XDC_R_0_146 VGND VNB vpwr_R_146 vpwr_R_146 sky130_fd_sc_hd__decap_12
XDC_R_1_146 VGND VNB vpwr_R_146 vpwr_R_146 sky130_fd_sc_hd__decap_12
XDC_R_2_146 VGND VNB vpwr_R_146 vpwr_R_146 sky130_fd_sc_hd__decap_12
XDC_R_0_147 VGND VNB vpwr_R_147 vpwr_R_147 sky130_fd_sc_hd__decap_12
XDC_R_1_147 VGND VNB vpwr_R_147 vpwr_R_147 sky130_fd_sc_hd__decap_12
XDC_R_2_147 VGND VNB vpwr_R_147 vpwr_R_147 sky130_fd_sc_hd__decap_12
XDC_R_0_148 VGND VNB vpwr_R_148 vpwr_R_148 sky130_fd_sc_hd__decap_12
XDC_R_1_148 VGND VNB vpwr_R_148 vpwr_R_148 sky130_fd_sc_hd__decap_12
XDC_R_2_148 VGND VNB vpwr_R_148 vpwr_R_148 sky130_fd_sc_hd__decap_12
XDC_R_0_149 VGND VNB vpwr_R_149 vpwr_R_149 sky130_fd_sc_hd__decap_12
XDC_R_1_149 VGND VNB vpwr_R_149 vpwr_R_149 sky130_fd_sc_hd__decap_12
XDC_R_2_149 VGND VNB vpwr_R_149 vpwr_R_149 sky130_fd_sc_hd__decap_12
XDC_R_0_150 VGND VNB vpwr_R_150 vpwr_R_150 sky130_fd_sc_hd__decap_12
XDC_R_1_150 VGND VNB vpwr_R_150 vpwr_R_150 sky130_fd_sc_hd__decap_12
XDC_R_2_150 VGND VNB vpwr_R_150 vpwr_R_150 sky130_fd_sc_hd__decap_12
XDC_R_0_151 VGND VNB vpwr_R_151 vpwr_R_151 sky130_fd_sc_hd__decap_12
XDC_R_1_151 VGND VNB vpwr_R_151 vpwr_R_151 sky130_fd_sc_hd__decap_12
XDC_R_2_151 VGND VNB vpwr_R_151 vpwr_R_151 sky130_fd_sc_hd__decap_12
XDC_R_0_152 VGND VNB vpwr_R_152 vpwr_R_152 sky130_fd_sc_hd__decap_12
XDC_R_1_152 VGND VNB vpwr_R_152 vpwr_R_152 sky130_fd_sc_hd__decap_12
XDC_R_2_152 VGND VNB vpwr_R_152 vpwr_R_152 sky130_fd_sc_hd__decap_12
XDC_R_0_153 VGND VNB vpwr_R_153 vpwr_R_153 sky130_fd_sc_hd__decap_12
XDC_R_1_153 VGND VNB vpwr_R_153 vpwr_R_153 sky130_fd_sc_hd__decap_12
XDC_R_2_153 VGND VNB vpwr_R_153 vpwr_R_153 sky130_fd_sc_hd__decap_12
XDC_R_0_154 VGND VNB vpwr_R_154 vpwr_R_154 sky130_fd_sc_hd__decap_12
XDC_R_1_154 VGND VNB vpwr_R_154 vpwr_R_154 sky130_fd_sc_hd__decap_12
XDC_R_2_154 VGND VNB vpwr_R_154 vpwr_R_154 sky130_fd_sc_hd__decap_12
XDC_R_0_155 VGND VNB vpwr_R_155 vpwr_R_155 sky130_fd_sc_hd__decap_12
XDC_R_1_155 VGND VNB vpwr_R_155 vpwr_R_155 sky130_fd_sc_hd__decap_12
XDC_R_2_155 VGND VNB vpwr_R_155 vpwr_R_155 sky130_fd_sc_hd__decap_12
XDC_R_0_156 VGND VNB vpwr_R_156 vpwr_R_156 sky130_fd_sc_hd__decap_12
XDC_R_1_156 VGND VNB vpwr_R_156 vpwr_R_156 sky130_fd_sc_hd__decap_12
XDC_R_2_156 VGND VNB vpwr_R_156 vpwr_R_156 sky130_fd_sc_hd__decap_12
XDC_R_0_157 VGND VNB vpwr_R_157 vpwr_R_157 sky130_fd_sc_hd__decap_12
XDC_R_1_157 VGND VNB vpwr_R_157 vpwr_R_157 sky130_fd_sc_hd__decap_12
XDC_R_2_157 VGND VNB vpwr_R_157 vpwr_R_157 sky130_fd_sc_hd__decap_12
XDC_R_0_158 VGND VNB vpwr_R_158 vpwr_R_158 sky130_fd_sc_hd__decap_12
XDC_R_1_158 VGND VNB vpwr_R_158 vpwr_R_158 sky130_fd_sc_hd__decap_12
XDC_R_2_158 VGND VNB vpwr_R_158 vpwr_R_158 sky130_fd_sc_hd__decap_12
XDC_R_0_159 VGND VNB vpwr_R_159 vpwr_R_159 sky130_fd_sc_hd__decap_12
XDC_R_1_159 VGND VNB vpwr_R_159 vpwr_R_159 sky130_fd_sc_hd__decap_12
XDC_R_2_159 VGND VNB vpwr_R_159 vpwr_R_159 sky130_fd_sc_hd__decap_12
XDC_R_0_160 VGND VNB vpwr_R_160 vpwr_R_160 sky130_fd_sc_hd__decap_12
XDC_R_1_160 VGND VNB vpwr_R_160 vpwr_R_160 sky130_fd_sc_hd__decap_12
XDC_R_2_160 VGND VNB vpwr_R_160 vpwr_R_160 sky130_fd_sc_hd__decap_12
XDC_R_0_161 VGND VNB vpwr_R_161 vpwr_R_161 sky130_fd_sc_hd__decap_12
XDC_R_1_161 VGND VNB vpwr_R_161 vpwr_R_161 sky130_fd_sc_hd__decap_12
XDC_R_2_161 VGND VNB vpwr_R_161 vpwr_R_161 sky130_fd_sc_hd__decap_12
XDC_R_0_162 VGND VNB vpwr_R_162 vpwr_R_162 sky130_fd_sc_hd__decap_12
XDC_R_1_162 VGND VNB vpwr_R_162 vpwr_R_162 sky130_fd_sc_hd__decap_12
XDC_R_2_162 VGND VNB vpwr_R_162 vpwr_R_162 sky130_fd_sc_hd__decap_12
XDC_R_0_163 VGND VNB vpwr_R_163 vpwr_R_163 sky130_fd_sc_hd__decap_12
XDC_R_1_163 VGND VNB vpwr_R_163 vpwr_R_163 sky130_fd_sc_hd__decap_12
XDC_R_2_163 VGND VNB vpwr_R_163 vpwr_R_163 sky130_fd_sc_hd__decap_12
XDC_R_0_164 VGND VNB vpwr_R_164 vpwr_R_164 sky130_fd_sc_hd__decap_12
XDC_R_1_164 VGND VNB vpwr_R_164 vpwr_R_164 sky130_fd_sc_hd__decap_12
XDC_R_2_164 VGND VNB vpwr_R_164 vpwr_R_164 sky130_fd_sc_hd__decap_12
XDC_R_0_165 VGND VNB vpwr_R_165 vpwr_R_165 sky130_fd_sc_hd__decap_12
XDC_R_1_165 VGND VNB vpwr_R_165 vpwr_R_165 sky130_fd_sc_hd__decap_12
XDC_R_2_165 VGND VNB vpwr_R_165 vpwr_R_165 sky130_fd_sc_hd__decap_12
XDC_R_0_166 VGND VNB vpwr_R_166 vpwr_R_166 sky130_fd_sc_hd__decap_12
XDC_R_1_166 VGND VNB vpwr_R_166 vpwr_R_166 sky130_fd_sc_hd__decap_12
XDC_R_2_166 VGND VNB vpwr_R_166 vpwr_R_166 sky130_fd_sc_hd__decap_12
XDC_R_0_167 VGND VNB vpwr_R_167 vpwr_R_167 sky130_fd_sc_hd__decap_12
XDC_R_1_167 VGND VNB vpwr_R_167 vpwr_R_167 sky130_fd_sc_hd__decap_12
XDC_R_2_167 VGND VNB vpwr_R_167 vpwr_R_167 sky130_fd_sc_hd__decap_12
XDC_R_0_168 VGND VNB vpwr_R_168 vpwr_R_168 sky130_fd_sc_hd__decap_12
XDC_R_1_168 VGND VNB vpwr_R_168 vpwr_R_168 sky130_fd_sc_hd__decap_12
XDC_R_2_168 VGND VNB vpwr_R_168 vpwr_R_168 sky130_fd_sc_hd__decap_12
XDC_R_0_169 VGND VNB vpwr_R_169 vpwr_R_169 sky130_fd_sc_hd__decap_12
XDC_R_1_169 VGND VNB vpwr_R_169 vpwr_R_169 sky130_fd_sc_hd__decap_12
XDC_R_2_169 VGND VNB vpwr_R_169 vpwr_R_169 sky130_fd_sc_hd__decap_12
XDC_R_0_170 VGND VNB vpwr_R_170 vpwr_R_170 sky130_fd_sc_hd__decap_12
XDC_R_1_170 VGND VNB vpwr_R_170 vpwr_R_170 sky130_fd_sc_hd__decap_12
XDC_R_2_170 VGND VNB vpwr_R_170 vpwr_R_170 sky130_fd_sc_hd__decap_12
XDC_R_0_171 VGND VNB vpwr_R_171 vpwr_R_171 sky130_fd_sc_hd__decap_12
XDC_R_1_171 VGND VNB vpwr_R_171 vpwr_R_171 sky130_fd_sc_hd__decap_12
XDC_R_2_171 VGND VNB vpwr_R_171 vpwr_R_171 sky130_fd_sc_hd__decap_12
XDC_R_0_172 VGND VNB vpwr_R_172 vpwr_R_172 sky130_fd_sc_hd__decap_12
XDC_R_1_172 VGND VNB vpwr_R_172 vpwr_R_172 sky130_fd_sc_hd__decap_12
XDC_R_2_172 VGND VNB vpwr_R_172 vpwr_R_172 sky130_fd_sc_hd__decap_12
XDC_R_0_173 VGND VNB vpwr_R_173 vpwr_R_173 sky130_fd_sc_hd__decap_12
XDC_R_1_173 VGND VNB vpwr_R_173 vpwr_R_173 sky130_fd_sc_hd__decap_12
XDC_R_2_173 VGND VNB vpwr_R_173 vpwr_R_173 sky130_fd_sc_hd__decap_12
XDC_R_0_174 VGND VNB vpwr_R_174 vpwr_R_174 sky130_fd_sc_hd__decap_12
XDC_R_1_174 VGND VNB vpwr_R_174 vpwr_R_174 sky130_fd_sc_hd__decap_12
XDC_R_2_174 VGND VNB vpwr_R_174 vpwr_R_174 sky130_fd_sc_hd__decap_12
XDC_R_0_175 VGND VNB vpwr_R_175 vpwr_R_175 sky130_fd_sc_hd__decap_12
XDC_R_1_175 VGND VNB vpwr_R_175 vpwr_R_175 sky130_fd_sc_hd__decap_12
XDC_R_2_175 VGND VNB vpwr_R_175 vpwr_R_175 sky130_fd_sc_hd__decap_12
XDC_R_0_176 VGND VNB vpwr_R_176 vpwr_R_176 sky130_fd_sc_hd__decap_12
XDC_R_1_176 VGND VNB vpwr_R_176 vpwr_R_176 sky130_fd_sc_hd__decap_12
XDC_R_2_176 VGND VNB vpwr_R_176 vpwr_R_176 sky130_fd_sc_hd__decap_12
XDC_R_0_177 VGND VNB vpwr_R_177 vpwr_R_177 sky130_fd_sc_hd__decap_12
XDC_R_1_177 VGND VNB vpwr_R_177 vpwr_R_177 sky130_fd_sc_hd__decap_12
XDC_R_2_177 VGND VNB vpwr_R_177 vpwr_R_177 sky130_fd_sc_hd__decap_12
XDC_R_0_178 VGND VNB vpwr_R_178 vpwr_R_178 sky130_fd_sc_hd__decap_12
XDC_R_1_178 VGND VNB vpwr_R_178 vpwr_R_178 sky130_fd_sc_hd__decap_12
XDC_R_2_178 VGND VNB vpwr_R_178 vpwr_R_178 sky130_fd_sc_hd__decap_12
XDC_R_0_179 VGND VNB vpwr_R_179 vpwr_R_179 sky130_fd_sc_hd__decap_12
XDC_R_1_179 VGND VNB vpwr_R_179 vpwr_R_179 sky130_fd_sc_hd__decap_12
XDC_R_2_179 VGND VNB vpwr_R_179 vpwr_R_179 sky130_fd_sc_hd__decap_12
XDC_R_0_180 VGND VNB vpwr_R_180 vpwr_R_180 sky130_fd_sc_hd__decap_12
XDC_R_1_180 VGND VNB vpwr_R_180 vpwr_R_180 sky130_fd_sc_hd__decap_12
XDC_R_2_180 VGND VNB vpwr_R_180 vpwr_R_180 sky130_fd_sc_hd__decap_12
XDC_R_0_181 VGND VNB vpwr_R_181 vpwr_R_181 sky130_fd_sc_hd__decap_12
XDC_R_1_181 VGND VNB vpwr_R_181 vpwr_R_181 sky130_fd_sc_hd__decap_12
XDC_R_2_181 VGND VNB vpwr_R_181 vpwr_R_181 sky130_fd_sc_hd__decap_12
XDC_R_0_182 VGND VNB vpwr_R_182 vpwr_R_182 sky130_fd_sc_hd__decap_12
XDC_R_1_182 VGND VNB vpwr_R_182 vpwr_R_182 sky130_fd_sc_hd__decap_12
XDC_R_2_182 VGND VNB vpwr_R_182 vpwr_R_182 sky130_fd_sc_hd__decap_12
XDC_R_0_183 VGND VNB vpwr_R_183 vpwr_R_183 sky130_fd_sc_hd__decap_12
XDC_R_1_183 VGND VNB vpwr_R_183 vpwr_R_183 sky130_fd_sc_hd__decap_12
XDC_R_2_183 VGND VNB vpwr_R_183 vpwr_R_183 sky130_fd_sc_hd__decap_12
XDC_R_0_184 VGND VNB vpwr_R_184 vpwr_R_184 sky130_fd_sc_hd__decap_12
XDC_R_1_184 VGND VNB vpwr_R_184 vpwr_R_184 sky130_fd_sc_hd__decap_12
XDC_R_2_184 VGND VNB vpwr_R_184 vpwr_R_184 sky130_fd_sc_hd__decap_12
XDC_R_0_185 VGND VNB vpwr_R_185 vpwr_R_185 sky130_fd_sc_hd__decap_12
XDC_R_1_185 VGND VNB vpwr_R_185 vpwr_R_185 sky130_fd_sc_hd__decap_12
XDC_R_2_185 VGND VNB vpwr_R_185 vpwr_R_185 sky130_fd_sc_hd__decap_12
XDC_R_0_186 VGND VNB vpwr_R_186 vpwr_R_186 sky130_fd_sc_hd__decap_12
XDC_R_1_186 VGND VNB vpwr_R_186 vpwr_R_186 sky130_fd_sc_hd__decap_12
XDC_R_2_186 VGND VNB vpwr_R_186 vpwr_R_186 sky130_fd_sc_hd__decap_12
XDC_R_0_187 VGND VNB vpwr_R_187 vpwr_R_187 sky130_fd_sc_hd__decap_12
XDC_R_1_187 VGND VNB vpwr_R_187 vpwr_R_187 sky130_fd_sc_hd__decap_12
XDC_R_2_187 VGND VNB vpwr_R_187 vpwr_R_187 sky130_fd_sc_hd__decap_12
XDC_R_0_188 VGND VNB vpwr_R_188 vpwr_R_188 sky130_fd_sc_hd__decap_12
XDC_R_1_188 VGND VNB vpwr_R_188 vpwr_R_188 sky130_fd_sc_hd__decap_12
XDC_R_2_188 VGND VNB vpwr_R_188 vpwr_R_188 sky130_fd_sc_hd__decap_12
XDC_R_0_189 VGND VNB vpwr_R_189 vpwr_R_189 sky130_fd_sc_hd__decap_12
XDC_R_1_189 VGND VNB vpwr_R_189 vpwr_R_189 sky130_fd_sc_hd__decap_12
XDC_R_2_189 VGND VNB vpwr_R_189 vpwr_R_189 sky130_fd_sc_hd__decap_12
XDC_R_0_190 VGND VNB vpwr_R_190 vpwr_R_190 sky130_fd_sc_hd__decap_12
XDC_R_1_190 VGND VNB vpwr_R_190 vpwr_R_190 sky130_fd_sc_hd__decap_12
XDC_R_2_190 VGND VNB vpwr_R_190 vpwr_R_190 sky130_fd_sc_hd__decap_12
XDC_R_0_191 VGND VNB vpwr_R_191 vpwr_R_191 sky130_fd_sc_hd__decap_12
XDC_R_1_191 VGND VNB vpwr_R_191 vpwr_R_191 sky130_fd_sc_hd__decap_12
XDC_R_2_191 VGND VNB vpwr_R_191 vpwr_R_191 sky130_fd_sc_hd__decap_12
XDC_R_0_192 VGND VNB vpwr_R_192 vpwr_R_192 sky130_fd_sc_hd__decap_12
XDC_R_1_192 VGND VNB vpwr_R_192 vpwr_R_192 sky130_fd_sc_hd__decap_12
XDC_R_2_192 VGND VNB vpwr_R_192 vpwr_R_192 sky130_fd_sc_hd__decap_12
XDC_R_0_193 VGND VNB vpwr_R_193 vpwr_R_193 sky130_fd_sc_hd__decap_12
XDC_R_1_193 VGND VNB vpwr_R_193 vpwr_R_193 sky130_fd_sc_hd__decap_12
XDC_R_2_193 VGND VNB vpwr_R_193 vpwr_R_193 sky130_fd_sc_hd__decap_12
XDC_R_0_194 VGND VNB vpwr_R_194 vpwr_R_194 sky130_fd_sc_hd__decap_12
XDC_R_1_194 VGND VNB vpwr_R_194 vpwr_R_194 sky130_fd_sc_hd__decap_12
XDC_R_2_194 VGND VNB vpwr_R_194 vpwr_R_194 sky130_fd_sc_hd__decap_12
XDC_R_0_195 VGND VNB vpwr_R_195 vpwr_R_195 sky130_fd_sc_hd__decap_12
XDC_R_1_195 VGND VNB vpwr_R_195 vpwr_R_195 sky130_fd_sc_hd__decap_12
XDC_R_2_195 VGND VNB vpwr_R_195 vpwr_R_195 sky130_fd_sc_hd__decap_12
XDC_R_0_196 VGND VNB vpwr_R_196 vpwr_R_196 sky130_fd_sc_hd__decap_12
XDC_R_1_196 VGND VNB vpwr_R_196 vpwr_R_196 sky130_fd_sc_hd__decap_12
XDC_R_2_196 VGND VNB vpwr_R_196 vpwr_R_196 sky130_fd_sc_hd__decap_12
XDC_R_0_197 VGND VNB vpwr_R_197 vpwr_R_197 sky130_fd_sc_hd__decap_12
XDC_R_1_197 VGND VNB vpwr_R_197 vpwr_R_197 sky130_fd_sc_hd__decap_12
XDC_R_2_197 VGND VNB vpwr_R_197 vpwr_R_197 sky130_fd_sc_hd__decap_12
XDC_R_0_198 VGND VNB vpwr_R_198 vpwr_R_198 sky130_fd_sc_hd__decap_12
XDC_R_1_198 VGND VNB vpwr_R_198 vpwr_R_198 sky130_fd_sc_hd__decap_12
XDC_R_2_198 VGND VNB vpwr_R_198 vpwr_R_198 sky130_fd_sc_hd__decap_12
XDC_R_0_199 VGND VNB vpwr_R_199 vpwr_R_199 sky130_fd_sc_hd__decap_12
XDC_R_1_199 VGND VNB vpwr_R_199 vpwr_R_199 sky130_fd_sc_hd__decap_12
XDC_R_2_199 VGND VNB vpwr_R_199 vpwr_R_199 sky130_fd_sc_hd__decap_12
XDC_R_0_200 VGND VNB vpwr_R_200 vpwr_R_200 sky130_fd_sc_hd__decap_12
XDC_R_1_200 VGND VNB vpwr_R_200 vpwr_R_200 sky130_fd_sc_hd__decap_12
XDC_R_2_200 VGND VNB vpwr_R_200 vpwr_R_200 sky130_fd_sc_hd__decap_12
XDC_R_0_201 VGND VNB vpwr_R_201 vpwr_R_201 sky130_fd_sc_hd__decap_12
XDC_R_1_201 VGND VNB vpwr_R_201 vpwr_R_201 sky130_fd_sc_hd__decap_12
XDC_R_2_201 VGND VNB vpwr_R_201 vpwr_R_201 sky130_fd_sc_hd__decap_12
XDC_R_0_202 VGND VNB vpwr_R_202 vpwr_R_202 sky130_fd_sc_hd__decap_12
XDC_R_1_202 VGND VNB vpwr_R_202 vpwr_R_202 sky130_fd_sc_hd__decap_12
XDC_R_2_202 VGND VNB vpwr_R_202 vpwr_R_202 sky130_fd_sc_hd__decap_12
XDC_R_0_203 VGND VNB vpwr_R_203 vpwr_R_203 sky130_fd_sc_hd__decap_12
XDC_R_1_203 VGND VNB vpwr_R_203 vpwr_R_203 sky130_fd_sc_hd__decap_12
XDC_R_2_203 VGND VNB vpwr_R_203 vpwr_R_203 sky130_fd_sc_hd__decap_12
XDC_R_0_204 VGND VNB vpwr_R_204 vpwr_R_204 sky130_fd_sc_hd__decap_12
XDC_R_1_204 VGND VNB vpwr_R_204 vpwr_R_204 sky130_fd_sc_hd__decap_12
XDC_R_2_204 VGND VNB vpwr_R_204 vpwr_R_204 sky130_fd_sc_hd__decap_12
XDC_R_0_205 VGND VNB vpwr_R_205 vpwr_R_205 sky130_fd_sc_hd__decap_12
XDC_R_1_205 VGND VNB vpwr_R_205 vpwr_R_205 sky130_fd_sc_hd__decap_12
XDC_R_2_205 VGND VNB vpwr_R_205 vpwr_R_205 sky130_fd_sc_hd__decap_12
XDC_R_0_206 VGND VNB vpwr_R_206 vpwr_R_206 sky130_fd_sc_hd__decap_12
XDC_R_1_206 VGND VNB vpwr_R_206 vpwr_R_206 sky130_fd_sc_hd__decap_12
XDC_R_2_206 VGND VNB vpwr_R_206 vpwr_R_206 sky130_fd_sc_hd__decap_12
XDC_R_0_207 VGND VNB vpwr_R_207 vpwr_R_207 sky130_fd_sc_hd__decap_12
XDC_R_1_207 VGND VNB vpwr_R_207 vpwr_R_207 sky130_fd_sc_hd__decap_12
XDC_R_2_207 VGND VNB vpwr_R_207 vpwr_R_207 sky130_fd_sc_hd__decap_12
XDC_R_0_208 VGND VNB vpwr_R_208 vpwr_R_208 sky130_fd_sc_hd__decap_12
XDC_R_1_208 VGND VNB vpwr_R_208 vpwr_R_208 sky130_fd_sc_hd__decap_12
XDC_R_2_208 VGND VNB vpwr_R_208 vpwr_R_208 sky130_fd_sc_hd__decap_12
XDC_R_0_209 VGND VNB vpwr_R_209 vpwr_R_209 sky130_fd_sc_hd__decap_12
XDC_R_1_209 VGND VNB vpwr_R_209 vpwr_R_209 sky130_fd_sc_hd__decap_12
XDC_R_2_209 VGND VNB vpwr_R_209 vpwr_R_209 sky130_fd_sc_hd__decap_12
XDC_R_0_210 VGND VNB vpwr_R_210 vpwr_R_210 sky130_fd_sc_hd__decap_12
XDC_R_1_210 VGND VNB vpwr_R_210 vpwr_R_210 sky130_fd_sc_hd__decap_12
XDC_R_2_210 VGND VNB vpwr_R_210 vpwr_R_210 sky130_fd_sc_hd__decap_12
XDC_R_0_211 VGND VNB vpwr_R_211 vpwr_R_211 sky130_fd_sc_hd__decap_12
XDC_R_1_211 VGND VNB vpwr_R_211 vpwr_R_211 sky130_fd_sc_hd__decap_12
XDC_R_2_211 VGND VNB vpwr_R_211 vpwr_R_211 sky130_fd_sc_hd__decap_12
XDC_R_0_212 VGND VNB vpwr_R_212 vpwr_R_212 sky130_fd_sc_hd__decap_12
XDC_R_1_212 VGND VNB vpwr_R_212 vpwr_R_212 sky130_fd_sc_hd__decap_12
XDC_R_2_212 VGND VNB vpwr_R_212 vpwr_R_212 sky130_fd_sc_hd__decap_12
XDC_R_0_213 VGND VNB vpwr_R_213 vpwr_R_213 sky130_fd_sc_hd__decap_12
XDC_R_1_213 VGND VNB vpwr_R_213 vpwr_R_213 sky130_fd_sc_hd__decap_12
XDC_R_2_213 VGND VNB vpwr_R_213 vpwr_R_213 sky130_fd_sc_hd__decap_12
XDC_R_0_214 VGND VNB vpwr_R_214 vpwr_R_214 sky130_fd_sc_hd__decap_12
XDC_R_1_214 VGND VNB vpwr_R_214 vpwr_R_214 sky130_fd_sc_hd__decap_12
XDC_R_2_214 VGND VNB vpwr_R_214 vpwr_R_214 sky130_fd_sc_hd__decap_12
XDC_R_0_215 VGND VNB vpwr_R_215 vpwr_R_215 sky130_fd_sc_hd__decap_12
XDC_R_1_215 VGND VNB vpwr_R_215 vpwr_R_215 sky130_fd_sc_hd__decap_12
XDC_R_2_215 VGND VNB vpwr_R_215 vpwr_R_215 sky130_fd_sc_hd__decap_12
XDC_R_0_216 VGND VNB vpwr_R_216 vpwr_R_216 sky130_fd_sc_hd__decap_12
XDC_R_1_216 VGND VNB vpwr_R_216 vpwr_R_216 sky130_fd_sc_hd__decap_12
XDC_R_2_216 VGND VNB vpwr_R_216 vpwr_R_216 sky130_fd_sc_hd__decap_12
XDC_R_0_217 VGND VNB vpwr_R_217 vpwr_R_217 sky130_fd_sc_hd__decap_12
XDC_R_1_217 VGND VNB vpwr_R_217 vpwr_R_217 sky130_fd_sc_hd__decap_12
XDC_R_2_217 VGND VNB vpwr_R_217 vpwr_R_217 sky130_fd_sc_hd__decap_12
XDC_R_0_218 VGND VNB vpwr_R_218 vpwr_R_218 sky130_fd_sc_hd__decap_12
XDC_R_1_218 VGND VNB vpwr_R_218 vpwr_R_218 sky130_fd_sc_hd__decap_12
XDC_R_2_218 VGND VNB vpwr_R_218 vpwr_R_218 sky130_fd_sc_hd__decap_12
XDC_R_0_219 VGND VNB vpwr_R_219 vpwr_R_219 sky130_fd_sc_hd__decap_12
XDC_R_1_219 VGND VNB vpwr_R_219 vpwr_R_219 sky130_fd_sc_hd__decap_12
XDC_R_2_219 VGND VNB vpwr_R_219 vpwr_R_219 sky130_fd_sc_hd__decap_12
XDC_R_0_220 VGND VNB vpwr_R_220 vpwr_R_220 sky130_fd_sc_hd__decap_12
XDC_R_1_220 VGND VNB vpwr_R_220 vpwr_R_220 sky130_fd_sc_hd__decap_12
XDC_R_2_220 VGND VNB vpwr_R_220 vpwr_R_220 sky130_fd_sc_hd__decap_12
XDC_R_0_221 VGND VNB vpwr_R_221 vpwr_R_221 sky130_fd_sc_hd__decap_12
XDC_R_1_221 VGND VNB vpwr_R_221 vpwr_R_221 sky130_fd_sc_hd__decap_12
XDC_R_2_221 VGND VNB vpwr_R_221 vpwr_R_221 sky130_fd_sc_hd__decap_12
XDC_R_0_222 VGND VNB vpwr_R_222 vpwr_R_222 sky130_fd_sc_hd__decap_12
XDC_R_1_222 VGND VNB vpwr_R_222 vpwr_R_222 sky130_fd_sc_hd__decap_12
XDC_R_2_222 VGND VNB vpwr_R_222 vpwr_R_222 sky130_fd_sc_hd__decap_12
XDC_R_0_223 VGND VNB vpwr_R_223 vpwr_R_223 sky130_fd_sc_hd__decap_12
XDC_R_1_223 VGND VNB vpwr_R_223 vpwr_R_223 sky130_fd_sc_hd__decap_12
XDC_R_2_223 VGND VNB vpwr_R_223 vpwr_R_223 sky130_fd_sc_hd__decap_12
XDC_R_0_224 VGND VNB vpwr_R_224 vpwr_R_224 sky130_fd_sc_hd__decap_12
XDC_R_1_224 VGND VNB vpwr_R_224 vpwr_R_224 sky130_fd_sc_hd__decap_12
XDC_R_2_224 VGND VNB vpwr_R_224 vpwr_R_224 sky130_fd_sc_hd__decap_12
XDC_R_0_225 VGND VNB vpwr_R_225 vpwr_R_225 sky130_fd_sc_hd__decap_12
XDC_R_1_225 VGND VNB vpwr_R_225 vpwr_R_225 sky130_fd_sc_hd__decap_12
XDC_R_2_225 VGND VNB vpwr_R_225 vpwr_R_225 sky130_fd_sc_hd__decap_12
XDC_R_0_226 VGND VNB vpwr_R_226 vpwr_R_226 sky130_fd_sc_hd__decap_12
XDC_R_1_226 VGND VNB vpwr_R_226 vpwr_R_226 sky130_fd_sc_hd__decap_12
XDC_R_2_226 VGND VNB vpwr_R_226 vpwr_R_226 sky130_fd_sc_hd__decap_12
XDC_R_0_227 VGND VNB vpwr_R_227 vpwr_R_227 sky130_fd_sc_hd__decap_12
XDC_R_1_227 VGND VNB vpwr_R_227 vpwr_R_227 sky130_fd_sc_hd__decap_12
XDC_R_2_227 VGND VNB vpwr_R_227 vpwr_R_227 sky130_fd_sc_hd__decap_12
XDC_R_0_228 VGND VNB vpwr_R_228 vpwr_R_228 sky130_fd_sc_hd__decap_12
XDC_R_1_228 VGND VNB vpwr_R_228 vpwr_R_228 sky130_fd_sc_hd__decap_12
XDC_R_2_228 VGND VNB vpwr_R_228 vpwr_R_228 sky130_fd_sc_hd__decap_12
XDC_R_0_229 VGND VNB vpwr_R_229 vpwr_R_229 sky130_fd_sc_hd__decap_12
XDC_R_1_229 VGND VNB vpwr_R_229 vpwr_R_229 sky130_fd_sc_hd__decap_12
XDC_R_2_229 VGND VNB vpwr_R_229 vpwr_R_229 sky130_fd_sc_hd__decap_12
XDC_R_0_230 VGND VNB vpwr_R_230 vpwr_R_230 sky130_fd_sc_hd__decap_12
XDC_R_1_230 VGND VNB vpwr_R_230 vpwr_R_230 sky130_fd_sc_hd__decap_12
XDC_R_2_230 VGND VNB vpwr_R_230 vpwr_R_230 sky130_fd_sc_hd__decap_12
XDC_R_0_231 VGND VNB vpwr_R_231 vpwr_R_231 sky130_fd_sc_hd__decap_12
XDC_R_1_231 VGND VNB vpwr_R_231 vpwr_R_231 sky130_fd_sc_hd__decap_12
XDC_R_2_231 VGND VNB vpwr_R_231 vpwr_R_231 sky130_fd_sc_hd__decap_12
XDC_R_0_232 VGND VNB vpwr_R_232 vpwr_R_232 sky130_fd_sc_hd__decap_12
XDC_R_1_232 VGND VNB vpwr_R_232 vpwr_R_232 sky130_fd_sc_hd__decap_12
XDC_R_2_232 VGND VNB vpwr_R_232 vpwr_R_232 sky130_fd_sc_hd__decap_12
XDC_R_0_233 VGND VNB vpwr_R_233 vpwr_R_233 sky130_fd_sc_hd__decap_12
XDC_R_1_233 VGND VNB vpwr_R_233 vpwr_R_233 sky130_fd_sc_hd__decap_12
XDC_R_2_233 VGND VNB vpwr_R_233 vpwr_R_233 sky130_fd_sc_hd__decap_12
XDC_R_0_234 VGND VNB vpwr_R_234 vpwr_R_234 sky130_fd_sc_hd__decap_12
XDC_R_1_234 VGND VNB vpwr_R_234 vpwr_R_234 sky130_fd_sc_hd__decap_12
XDC_R_2_234 VGND VNB vpwr_R_234 vpwr_R_234 sky130_fd_sc_hd__decap_12
XDC_R_0_235 VGND VNB vpwr_R_235 vpwr_R_235 sky130_fd_sc_hd__decap_12
XDC_R_1_235 VGND VNB vpwr_R_235 vpwr_R_235 sky130_fd_sc_hd__decap_12
XDC_R_2_235 VGND VNB vpwr_R_235 vpwr_R_235 sky130_fd_sc_hd__decap_12
XDC_R_0_236 VGND VNB vpwr_R_236 vpwr_R_236 sky130_fd_sc_hd__decap_12
XDC_R_1_236 VGND VNB vpwr_R_236 vpwr_R_236 sky130_fd_sc_hd__decap_12
XDC_R_2_236 VGND VNB vpwr_R_236 vpwr_R_236 sky130_fd_sc_hd__decap_12
XDC_R_0_237 VGND VNB vpwr_R_237 vpwr_R_237 sky130_fd_sc_hd__decap_12
XDC_R_1_237 VGND VNB vpwr_R_237 vpwr_R_237 sky130_fd_sc_hd__decap_12
XDC_R_2_237 VGND VNB vpwr_R_237 vpwr_R_237 sky130_fd_sc_hd__decap_12
XDC_R_0_238 VGND VNB vpwr_R_238 vpwr_R_238 sky130_fd_sc_hd__decap_12
XDC_R_1_238 VGND VNB vpwr_R_238 vpwr_R_238 sky130_fd_sc_hd__decap_12
XDC_R_2_238 VGND VNB vpwr_R_238 vpwr_R_238 sky130_fd_sc_hd__decap_12
XDC_R_0_239 VGND VNB vpwr_R_239 vpwr_R_239 sky130_fd_sc_hd__decap_12
XDC_R_1_239 VGND VNB vpwr_R_239 vpwr_R_239 sky130_fd_sc_hd__decap_12
XDC_R_2_239 VGND VNB vpwr_R_239 vpwr_R_239 sky130_fd_sc_hd__decap_12
XDC_R_0_240 VGND VNB vpwr_R_240 vpwr_R_240 sky130_fd_sc_hd__decap_12
XDC_R_1_240 VGND VNB vpwr_R_240 vpwr_R_240 sky130_fd_sc_hd__decap_12
XDC_R_2_240 VGND VNB vpwr_R_240 vpwr_R_240 sky130_fd_sc_hd__decap_12
XDC_R_0_241 VGND VNB vpwr_R_241 vpwr_R_241 sky130_fd_sc_hd__decap_12
XDC_R_1_241 VGND VNB vpwr_R_241 vpwr_R_241 sky130_fd_sc_hd__decap_12
XDC_R_2_241 VGND VNB vpwr_R_241 vpwr_R_241 sky130_fd_sc_hd__decap_12
XDC_R_0_242 VGND VNB vpwr_R_242 vpwr_R_242 sky130_fd_sc_hd__decap_12
XDC_R_1_242 VGND VNB vpwr_R_242 vpwr_R_242 sky130_fd_sc_hd__decap_12
XDC_R_2_242 VGND VNB vpwr_R_242 vpwr_R_242 sky130_fd_sc_hd__decap_12
XDC_R_0_243 VGND VNB vpwr_R_243 vpwr_R_243 sky130_fd_sc_hd__decap_12
XDC_R_1_243 VGND VNB vpwr_R_243 vpwr_R_243 sky130_fd_sc_hd__decap_12
XDC_R_2_243 VGND VNB vpwr_R_243 vpwr_R_243 sky130_fd_sc_hd__decap_12
XDC_R_0_244 VGND VNB vpwr_R_244 vpwr_R_244 sky130_fd_sc_hd__decap_12
XDC_R_1_244 VGND VNB vpwr_R_244 vpwr_R_244 sky130_fd_sc_hd__decap_12
XDC_R_2_244 VGND VNB vpwr_R_244 vpwr_R_244 sky130_fd_sc_hd__decap_12
XDC_R_0_245 VGND VNB vpwr_R_245 vpwr_R_245 sky130_fd_sc_hd__decap_12
XDC_R_1_245 VGND VNB vpwr_R_245 vpwr_R_245 sky130_fd_sc_hd__decap_12
XDC_R_2_245 VGND VNB vpwr_R_245 vpwr_R_245 sky130_fd_sc_hd__decap_12
XDC_R_0_246 VGND VNB vpwr_R_246 vpwr_R_246 sky130_fd_sc_hd__decap_12
XDC_R_1_246 VGND VNB vpwr_R_246 vpwr_R_246 sky130_fd_sc_hd__decap_12
XDC_R_2_246 VGND VNB vpwr_R_246 vpwr_R_246 sky130_fd_sc_hd__decap_12
XDC_R_0_247 VGND VNB vpwr_R_247 vpwr_R_247 sky130_fd_sc_hd__decap_12
XDC_R_1_247 VGND VNB vpwr_R_247 vpwr_R_247 sky130_fd_sc_hd__decap_12
XDC_R_2_247 VGND VNB vpwr_R_247 vpwr_R_247 sky130_fd_sc_hd__decap_12
XDC_R_0_248 VGND VNB vpwr_R_248 vpwr_R_248 sky130_fd_sc_hd__decap_12
XDC_R_1_248 VGND VNB vpwr_R_248 vpwr_R_248 sky130_fd_sc_hd__decap_12
XDC_R_2_248 VGND VNB vpwr_R_248 vpwr_R_248 sky130_fd_sc_hd__decap_12
XDC_R_0_249 VGND VNB vpwr_R_249 vpwr_R_249 sky130_fd_sc_hd__decap_12
XDC_R_1_249 VGND VNB vpwr_R_249 vpwr_R_249 sky130_fd_sc_hd__decap_12
XDC_R_2_249 VGND VNB vpwr_R_249 vpwr_R_249 sky130_fd_sc_hd__decap_12
XDC_R_0_250 VGND VNB vpwr_R_250 vpwr_R_250 sky130_fd_sc_hd__decap_12
XDC_R_1_250 VGND VNB vpwr_R_250 vpwr_R_250 sky130_fd_sc_hd__decap_12
XDC_R_2_250 VGND VNB vpwr_R_250 vpwr_R_250 sky130_fd_sc_hd__decap_12
XDC_R_0_251 VGND VNB vpwr_R_251 vpwr_R_251 sky130_fd_sc_hd__decap_12
XDC_R_1_251 VGND VNB vpwr_R_251 vpwr_R_251 sky130_fd_sc_hd__decap_12
XDC_R_2_251 VGND VNB vpwr_R_251 vpwr_R_251 sky130_fd_sc_hd__decap_12
XDC_R_0_252 VGND VNB vpwr_R_252 vpwr_R_252 sky130_fd_sc_hd__decap_12
XDC_R_1_252 VGND VNB vpwr_R_252 vpwr_R_252 sky130_fd_sc_hd__decap_12
XDC_R_2_252 VGND VNB vpwr_R_252 vpwr_R_252 sky130_fd_sc_hd__decap_12
XDC_R_0_253 VGND VNB vpwr_R_253 vpwr_R_253 sky130_fd_sc_hd__decap_12
XDC_R_1_253 VGND VNB vpwr_R_253 vpwr_R_253 sky130_fd_sc_hd__decap_12
XDC_R_2_253 VGND VNB vpwr_R_253 vpwr_R_253 sky130_fd_sc_hd__decap_12
XDC_R_0_254 VGND VNB vpwr_R_254 vpwr_R_254 sky130_fd_sc_hd__decap_12
XDC_R_1_254 VGND VNB vpwr_R_254 vpwr_R_254 sky130_fd_sc_hd__decap_12
XDC_R_2_254 VGND VNB vpwr_R_254 vpwr_R_254 sky130_fd_sc_hd__decap_12
XDC_R_0_255 VGND VNB vpwr_R_255 vpwr_R_255 sky130_fd_sc_hd__decap_12
XDC_R_1_255 VGND VNB vpwr_R_255 vpwr_R_255 sky130_fd_sc_hd__decap_12
XDC_R_2_255 VGND VNB vpwr_R_255 vpwr_R_255 sky130_fd_sc_hd__decap_12
XDC_R_0_256 VGND VNB vpwr_R_256 vpwr_R_256 sky130_fd_sc_hd__decap_12
XDC_R_1_256 VGND VNB vpwr_R_256 vpwr_R_256 sky130_fd_sc_hd__decap_12
XDC_R_2_256 VGND VNB vpwr_R_256 vpwr_R_256 sky130_fd_sc_hd__decap_12
XDC_R_0_257 VGND VNB vpwr_R_257 vpwr_R_257 sky130_fd_sc_hd__decap_12
XDC_R_1_257 VGND VNB vpwr_R_257 vpwr_R_257 sky130_fd_sc_hd__decap_12
XDC_R_2_257 VGND VNB vpwr_R_257 vpwr_R_257 sky130_fd_sc_hd__decap_12
XDC_R_0_258 VGND VNB vpwr_R_258 vpwr_R_258 sky130_fd_sc_hd__decap_12
XDC_R_1_258 VGND VNB vpwr_R_258 vpwr_R_258 sky130_fd_sc_hd__decap_12
XDC_R_2_258 VGND VNB vpwr_R_258 vpwr_R_258 sky130_fd_sc_hd__decap_12
XDC_R_0_259 VGND VNB vpwr_R_259 vpwr_R_259 sky130_fd_sc_hd__decap_12
XDC_R_1_259 VGND VNB vpwr_R_259 vpwr_R_259 sky130_fd_sc_hd__decap_12
XDC_R_2_259 VGND VNB vpwr_R_259 vpwr_R_259 sky130_fd_sc_hd__decap_12
XDC_R_0_260 VGND VNB vpwr_R_260 vpwr_R_260 sky130_fd_sc_hd__decap_12
XDC_R_1_260 VGND VNB vpwr_R_260 vpwr_R_260 sky130_fd_sc_hd__decap_12
XDC_R_2_260 VGND VNB vpwr_R_260 vpwr_R_260 sky130_fd_sc_hd__decap_12
XDC_R_0_261 VGND VNB vpwr_R_261 vpwr_R_261 sky130_fd_sc_hd__decap_12
XDC_R_1_261 VGND VNB vpwr_R_261 vpwr_R_261 sky130_fd_sc_hd__decap_12
XDC_R_2_261 VGND VNB vpwr_R_261 vpwr_R_261 sky130_fd_sc_hd__decap_12
XDC_R_0_262 VGND VNB vpwr_R_262 vpwr_R_262 sky130_fd_sc_hd__decap_12
XDC_R_1_262 VGND VNB vpwr_R_262 vpwr_R_262 sky130_fd_sc_hd__decap_12
XDC_R_2_262 VGND VNB vpwr_R_262 vpwr_R_262 sky130_fd_sc_hd__decap_12
XDC_R_0_263 VGND VNB vpwr_R_263 vpwr_R_263 sky130_fd_sc_hd__decap_12
XDC_R_1_263 VGND VNB vpwr_R_263 vpwr_R_263 sky130_fd_sc_hd__decap_12
XDC_R_2_263 VGND VNB vpwr_R_263 vpwr_R_263 sky130_fd_sc_hd__decap_12
XDC_R_0_264 VGND VNB vpwr_R_264 vpwr_R_264 sky130_fd_sc_hd__decap_12
XDC_R_1_264 VGND VNB vpwr_R_264 vpwr_R_264 sky130_fd_sc_hd__decap_12
XDC_R_2_264 VGND VNB vpwr_R_264 vpwr_R_264 sky130_fd_sc_hd__decap_12
XDC_R_0_265 VGND VNB vpwr_R_265 vpwr_R_265 sky130_fd_sc_hd__decap_12
XDC_R_1_265 VGND VNB vpwr_R_265 vpwr_R_265 sky130_fd_sc_hd__decap_12
XDC_R_2_265 VGND VNB vpwr_R_265 vpwr_R_265 sky130_fd_sc_hd__decap_12
XDC_R_0_266 VGND VNB vpwr_R_266 vpwr_R_266 sky130_fd_sc_hd__decap_12
XDC_R_1_266 VGND VNB vpwr_R_266 vpwr_R_266 sky130_fd_sc_hd__decap_12
XDC_R_2_266 VGND VNB vpwr_R_266 vpwr_R_266 sky130_fd_sc_hd__decap_12
XDC_R_0_267 VGND VNB vpwr_R_267 vpwr_R_267 sky130_fd_sc_hd__decap_12
XDC_R_1_267 VGND VNB vpwr_R_267 vpwr_R_267 sky130_fd_sc_hd__decap_12
XDC_R_2_267 VGND VNB vpwr_R_267 vpwr_R_267 sky130_fd_sc_hd__decap_12
XDC_R_0_268 VGND VNB vpwr_R_268 vpwr_R_268 sky130_fd_sc_hd__decap_12
XDC_R_1_268 VGND VNB vpwr_R_268 vpwr_R_268 sky130_fd_sc_hd__decap_12
XDC_R_2_268 VGND VNB vpwr_R_268 vpwr_R_268 sky130_fd_sc_hd__decap_12
XDC_R_0_269 VGND VNB vpwr_R_269 vpwr_R_269 sky130_fd_sc_hd__decap_12
XDC_R_1_269 VGND VNB vpwr_R_269 vpwr_R_269 sky130_fd_sc_hd__decap_12
XDC_R_2_269 VGND VNB vpwr_R_269 vpwr_R_269 sky130_fd_sc_hd__decap_12
XDC_R_0_270 VGND VNB vpwr_R_270 vpwr_R_270 sky130_fd_sc_hd__decap_12
XDC_R_1_270 VGND VNB vpwr_R_270 vpwr_R_270 sky130_fd_sc_hd__decap_12
XDC_R_2_270 VGND VNB vpwr_R_270 vpwr_R_270 sky130_fd_sc_hd__decap_12
XDC_R_0_271 VGND VNB vpwr_R_271 vpwr_R_271 sky130_fd_sc_hd__decap_12
XDC_R_1_271 VGND VNB vpwr_R_271 vpwr_R_271 sky130_fd_sc_hd__decap_12
XDC_R_2_271 VGND VNB vpwr_R_271 vpwr_R_271 sky130_fd_sc_hd__decap_12
XDC_R_0_272 VGND VNB vpwr_R_272 vpwr_R_272 sky130_fd_sc_hd__decap_12
XDC_R_1_272 VGND VNB vpwr_R_272 vpwr_R_272 sky130_fd_sc_hd__decap_12
XDC_R_2_272 VGND VNB vpwr_R_272 vpwr_R_272 sky130_fd_sc_hd__decap_12
XDC_R_0_273 VGND VNB vpwr_R_273 vpwr_R_273 sky130_fd_sc_hd__decap_12
XDC_R_1_273 VGND VNB vpwr_R_273 vpwr_R_273 sky130_fd_sc_hd__decap_12
XDC_R_2_273 VGND VNB vpwr_R_273 vpwr_R_273 sky130_fd_sc_hd__decap_12
XDC_R_0_274 VGND VNB vpwr_R_274 vpwr_R_274 sky130_fd_sc_hd__decap_12
XDC_R_1_274 VGND VNB vpwr_R_274 vpwr_R_274 sky130_fd_sc_hd__decap_12
XDC_R_2_274 VGND VNB vpwr_R_274 vpwr_R_274 sky130_fd_sc_hd__decap_12
XDC_R_0_275 VGND VNB vpwr_R_275 vpwr_R_275 sky130_fd_sc_hd__decap_12
XDC_R_1_275 VGND VNB vpwr_R_275 vpwr_R_275 sky130_fd_sc_hd__decap_12
XDC_R_2_275 VGND VNB vpwr_R_275 vpwr_R_275 sky130_fd_sc_hd__decap_12
XDC_R_0_276 VGND VNB vpwr_R_276 vpwr_R_276 sky130_fd_sc_hd__decap_12
XDC_R_1_276 VGND VNB vpwr_R_276 vpwr_R_276 sky130_fd_sc_hd__decap_12
XDC_R_2_276 VGND VNB vpwr_R_276 vpwr_R_276 sky130_fd_sc_hd__decap_12
XDC_R_0_277 VGND VNB vpwr_R_277 vpwr_R_277 sky130_fd_sc_hd__decap_12
XDC_R_1_277 VGND VNB vpwr_R_277 vpwr_R_277 sky130_fd_sc_hd__decap_12
XDC_R_2_277 VGND VNB vpwr_R_277 vpwr_R_277 sky130_fd_sc_hd__decap_12
XDC_R_0_278 VGND VNB vpwr_R_278 vpwr_R_278 sky130_fd_sc_hd__decap_12
XDC_R_1_278 VGND VNB vpwr_R_278 vpwr_R_278 sky130_fd_sc_hd__decap_12
XDC_R_2_278 VGND VNB vpwr_R_278 vpwr_R_278 sky130_fd_sc_hd__decap_12
XDC_R_0_279 VGND VNB vpwr_R_279 vpwr_R_279 sky130_fd_sc_hd__decap_12
XDC_R_1_279 VGND VNB vpwr_R_279 vpwr_R_279 sky130_fd_sc_hd__decap_12
XDC_R_2_279 VGND VNB vpwr_R_279 vpwr_R_279 sky130_fd_sc_hd__decap_12
XDC_R_0_280 VGND VNB vpwr_R_280 vpwr_R_280 sky130_fd_sc_hd__decap_12
XDC_R_1_280 VGND VNB vpwr_R_280 vpwr_R_280 sky130_fd_sc_hd__decap_12
XDC_R_2_280 VGND VNB vpwr_R_280 vpwr_R_280 sky130_fd_sc_hd__decap_12
XDC_R_0_281 VGND VNB vpwr_R_281 vpwr_R_281 sky130_fd_sc_hd__decap_12
XDC_R_1_281 VGND VNB vpwr_R_281 vpwr_R_281 sky130_fd_sc_hd__decap_12
XDC_R_2_281 VGND VNB vpwr_R_281 vpwr_R_281 sky130_fd_sc_hd__decap_12
XDC_R_0_282 VGND VNB vpwr_R_282 vpwr_R_282 sky130_fd_sc_hd__decap_12
XDC_R_1_282 VGND VNB vpwr_R_282 vpwr_R_282 sky130_fd_sc_hd__decap_12
XDC_R_2_282 VGND VNB vpwr_R_282 vpwr_R_282 sky130_fd_sc_hd__decap_12
XDC_R_0_283 VGND VNB vpwr_R_283 vpwr_R_283 sky130_fd_sc_hd__decap_12
XDC_R_1_283 VGND VNB vpwr_R_283 vpwr_R_283 sky130_fd_sc_hd__decap_12
XDC_R_2_283 VGND VNB vpwr_R_283 vpwr_R_283 sky130_fd_sc_hd__decap_12
XDC_R_0_284 VGND VNB vpwr_R_284 vpwr_R_284 sky130_fd_sc_hd__decap_12
XDC_R_1_284 VGND VNB vpwr_R_284 vpwr_R_284 sky130_fd_sc_hd__decap_12
XDC_R_2_284 VGND VNB vpwr_R_284 vpwr_R_284 sky130_fd_sc_hd__decap_12
XDC_R_0_285 VGND VNB vpwr_R_285 vpwr_R_285 sky130_fd_sc_hd__decap_12
XDC_R_1_285 VGND VNB vpwr_R_285 vpwr_R_285 sky130_fd_sc_hd__decap_12
XDC_R_2_285 VGND VNB vpwr_R_285 vpwr_R_285 sky130_fd_sc_hd__decap_12
XDC_R_0_286 VGND VNB vpwr_R_286 vpwr_R_286 sky130_fd_sc_hd__decap_12
XDC_R_1_286 VGND VNB vpwr_R_286 vpwr_R_286 sky130_fd_sc_hd__decap_12
XDC_R_2_286 VGND VNB vpwr_R_286 vpwr_R_286 sky130_fd_sc_hd__decap_12
XDC_R_0_287 VGND VNB vpwr_R_287 vpwr_R_287 sky130_fd_sc_hd__decap_12
XDC_R_1_287 VGND VNB vpwr_R_287 vpwr_R_287 sky130_fd_sc_hd__decap_12
XDC_R_2_287 VGND VNB vpwr_R_287 vpwr_R_287 sky130_fd_sc_hd__decap_12
XDC_R_0_288 VGND VNB vpwr_R_288 vpwr_R_288 sky130_fd_sc_hd__decap_12
XDC_R_1_288 VGND VNB vpwr_R_288 vpwr_R_288 sky130_fd_sc_hd__decap_12
XDC_R_2_288 VGND VNB vpwr_R_288 vpwr_R_288 sky130_fd_sc_hd__decap_12
XDC_R_0_289 VGND VNB vpwr_R_289 vpwr_R_289 sky130_fd_sc_hd__decap_12
XDC_R_1_289 VGND VNB vpwr_R_289 vpwr_R_289 sky130_fd_sc_hd__decap_12
XDC_R_2_289 VGND VNB vpwr_R_289 vpwr_R_289 sky130_fd_sc_hd__decap_12
XDC_R_0_290 VGND VNB vpwr_R_290 vpwr_R_290 sky130_fd_sc_hd__decap_12
XDC_R_1_290 VGND VNB vpwr_R_290 vpwr_R_290 sky130_fd_sc_hd__decap_12
XDC_R_2_290 VGND VNB vpwr_R_290 vpwr_R_290 sky130_fd_sc_hd__decap_12
XDC_R_0_291 VGND VNB vpwr_R_291 vpwr_R_291 sky130_fd_sc_hd__decap_12
XDC_R_1_291 VGND VNB vpwr_R_291 vpwr_R_291 sky130_fd_sc_hd__decap_12
XDC_R_2_291 VGND VNB vpwr_R_291 vpwr_R_291 sky130_fd_sc_hd__decap_12
XDC_R_0_292 VGND VNB vpwr_R_292 vpwr_R_292 sky130_fd_sc_hd__decap_12
XDC_R_1_292 VGND VNB vpwr_R_292 vpwr_R_292 sky130_fd_sc_hd__decap_12
XDC_R_2_292 VGND VNB vpwr_R_292 vpwr_R_292 sky130_fd_sc_hd__decap_12
XDC_R_0_293 VGND VNB vpwr_R_293 vpwr_R_293 sky130_fd_sc_hd__decap_12
XDC_R_1_293 VGND VNB vpwr_R_293 vpwr_R_293 sky130_fd_sc_hd__decap_12
XDC_R_2_293 VGND VNB vpwr_R_293 vpwr_R_293 sky130_fd_sc_hd__decap_12
XDC_R_0_294 VGND VNB vpwr_R_294 vpwr_R_294 sky130_fd_sc_hd__decap_12
XDC_R_1_294 VGND VNB vpwr_R_294 vpwr_R_294 sky130_fd_sc_hd__decap_12
XDC_R_2_294 VGND VNB vpwr_R_294 vpwr_R_294 sky130_fd_sc_hd__decap_12
XDC_R_0_295 VGND VNB vpwr_R_295 vpwr_R_295 sky130_fd_sc_hd__decap_12
XDC_R_1_295 VGND VNB vpwr_R_295 vpwr_R_295 sky130_fd_sc_hd__decap_12
XDC_R_2_295 VGND VNB vpwr_R_295 vpwr_R_295 sky130_fd_sc_hd__decap_12
XDC_R_0_296 VGND VNB vpwr_R_296 vpwr_R_296 sky130_fd_sc_hd__decap_12
XDC_R_1_296 VGND VNB vpwr_R_296 vpwr_R_296 sky130_fd_sc_hd__decap_12
XDC_R_2_296 VGND VNB vpwr_R_296 vpwr_R_296 sky130_fd_sc_hd__decap_12
XDC_R_0_297 VGND VNB vpwr_R_297 vpwr_R_297 sky130_fd_sc_hd__decap_12
XDC_R_1_297 VGND VNB vpwr_R_297 vpwr_R_297 sky130_fd_sc_hd__decap_12
XDC_R_2_297 VGND VNB vpwr_R_297 vpwr_R_297 sky130_fd_sc_hd__decap_12
XDC_R_0_298 VGND VNB vpwr_R_298 vpwr_R_298 sky130_fd_sc_hd__decap_12
XDC_R_1_298 VGND VNB vpwr_R_298 vpwr_R_298 sky130_fd_sc_hd__decap_12
XDC_R_2_298 VGND VNB vpwr_R_298 vpwr_R_298 sky130_fd_sc_hd__decap_12
XDC_R_0_299 VGND VNB vpwr_R_299 vpwr_R_299 sky130_fd_sc_hd__decap_12
XDC_R_1_299 VGND VNB vpwr_R_299 vpwr_R_299 sky130_fd_sc_hd__decap_12
XDC_R_2_299 VGND VNB vpwr_R_299 vpwr_R_299 sky130_fd_sc_hd__decap_12
XDC_R_0_300 VGND VNB vpwr_R_300 vpwr_R_300 sky130_fd_sc_hd__decap_12
XDC_R_1_300 VGND VNB vpwr_R_300 vpwr_R_300 sky130_fd_sc_hd__decap_12
XDC_R_2_300 VGND VNB vpwr_R_300 vpwr_R_300 sky130_fd_sc_hd__decap_12
XDC_R_0_301 VGND VNB vpwr_R_301 vpwr_R_301 sky130_fd_sc_hd__decap_12
XDC_R_1_301 VGND VNB vpwr_R_301 vpwr_R_301 sky130_fd_sc_hd__decap_12
XDC_R_2_301 VGND VNB vpwr_R_301 vpwr_R_301 sky130_fd_sc_hd__decap_12
XDC_R_0_302 VGND VNB vpwr_R_302 vpwr_R_302 sky130_fd_sc_hd__decap_12
XDC_R_1_302 VGND VNB vpwr_R_302 vpwr_R_302 sky130_fd_sc_hd__decap_12
XDC_R_2_302 VGND VNB vpwr_R_302 vpwr_R_302 sky130_fd_sc_hd__decap_12
XDC_R_0_303 VGND VNB vpwr_R_303 vpwr_R_303 sky130_fd_sc_hd__decap_12
XDC_R_1_303 VGND VNB vpwr_R_303 vpwr_R_303 sky130_fd_sc_hd__decap_12
XDC_R_2_303 VGND VNB vpwr_R_303 vpwr_R_303 sky130_fd_sc_hd__decap_12
XDC_R_0_304 VGND VNB vpwr_R_304 vpwr_R_304 sky130_fd_sc_hd__decap_12
XDC_R_1_304 VGND VNB vpwr_R_304 vpwr_R_304 sky130_fd_sc_hd__decap_12
XDC_R_2_304 VGND VNB vpwr_R_304 vpwr_R_304 sky130_fd_sc_hd__decap_12
XDC_R_0_305 VGND VNB vpwr_R_305 vpwr_R_305 sky130_fd_sc_hd__decap_12
XDC_R_1_305 VGND VNB vpwr_R_305 vpwr_R_305 sky130_fd_sc_hd__decap_12
XDC_R_2_305 VGND VNB vpwr_R_305 vpwr_R_305 sky130_fd_sc_hd__decap_12
XDC_R_0_306 VGND VNB vpwr_R_306 vpwr_R_306 sky130_fd_sc_hd__decap_12
XDC_R_1_306 VGND VNB vpwr_R_306 vpwr_R_306 sky130_fd_sc_hd__decap_12
XDC_R_2_306 VGND VNB vpwr_R_306 vpwr_R_306 sky130_fd_sc_hd__decap_12
XDC_R_0_307 VGND VNB vpwr_R_307 vpwr_R_307 sky130_fd_sc_hd__decap_12
XDC_R_1_307 VGND VNB vpwr_R_307 vpwr_R_307 sky130_fd_sc_hd__decap_12
XDC_R_2_307 VGND VNB vpwr_R_307 vpwr_R_307 sky130_fd_sc_hd__decap_12
XDC_R_0_308 VGND VNB vpwr_R_308 vpwr_R_308 sky130_fd_sc_hd__decap_12
XDC_R_1_308 VGND VNB vpwr_R_308 vpwr_R_308 sky130_fd_sc_hd__decap_12
XDC_R_2_308 VGND VNB vpwr_R_308 vpwr_R_308 sky130_fd_sc_hd__decap_12
XDC_R_0_309 VGND VNB vpwr_R_309 vpwr_R_309 sky130_fd_sc_hd__decap_12
XDC_R_1_309 VGND VNB vpwr_R_309 vpwr_R_309 sky130_fd_sc_hd__decap_12
XDC_R_2_309 VGND VNB vpwr_R_309 vpwr_R_309 sky130_fd_sc_hd__decap_12
XDC_R_0_310 VGND VNB vpwr_R_310 vpwr_R_310 sky130_fd_sc_hd__decap_12
XDC_R_1_310 VGND VNB vpwr_R_310 vpwr_R_310 sky130_fd_sc_hd__decap_12
XDC_R_2_310 VGND VNB vpwr_R_310 vpwr_R_310 sky130_fd_sc_hd__decap_12
XDC_R_0_311 VGND VNB vpwr_R_311 vpwr_R_311 sky130_fd_sc_hd__decap_12
XDC_R_1_311 VGND VNB vpwr_R_311 vpwr_R_311 sky130_fd_sc_hd__decap_12
XDC_R_2_311 VGND VNB vpwr_R_311 vpwr_R_311 sky130_fd_sc_hd__decap_12
XDC_R_0_312 VGND VNB vpwr_R_312 vpwr_R_312 sky130_fd_sc_hd__decap_12
XDC_R_1_312 VGND VNB vpwr_R_312 vpwr_R_312 sky130_fd_sc_hd__decap_12
XDC_R_2_312 VGND VNB vpwr_R_312 vpwr_R_312 sky130_fd_sc_hd__decap_12
XDC_R_0_313 VGND VNB vpwr_R_313 vpwr_R_313 sky130_fd_sc_hd__decap_12
XDC_R_1_313 VGND VNB vpwr_R_313 vpwr_R_313 sky130_fd_sc_hd__decap_12
XDC_R_2_313 VGND VNB vpwr_R_313 vpwr_R_313 sky130_fd_sc_hd__decap_12
XDC_R_0_314 VGND VNB vpwr_R_314 vpwr_R_314 sky130_fd_sc_hd__decap_12
XDC_R_1_314 VGND VNB vpwr_R_314 vpwr_R_314 sky130_fd_sc_hd__decap_12
XDC_R_2_314 VGND VNB vpwr_R_314 vpwr_R_314 sky130_fd_sc_hd__decap_12
XDC_R_0_315 VGND VNB vpwr_R_315 vpwr_R_315 sky130_fd_sc_hd__decap_12
XDC_R_1_315 VGND VNB vpwr_R_315 vpwr_R_315 sky130_fd_sc_hd__decap_12
XDC_R_2_315 VGND VNB vpwr_R_315 vpwr_R_315 sky130_fd_sc_hd__decap_12
XDC_R_0_316 VGND VNB vpwr_R_316 vpwr_R_316 sky130_fd_sc_hd__decap_12
XDC_R_1_316 VGND VNB vpwr_R_316 vpwr_R_316 sky130_fd_sc_hd__decap_12
XDC_R_2_316 VGND VNB vpwr_R_316 vpwr_R_316 sky130_fd_sc_hd__decap_12
XDC_R_0_317 VGND VNB vpwr_R_317 vpwr_R_317 sky130_fd_sc_hd__decap_12
XDC_R_1_317 VGND VNB vpwr_R_317 vpwr_R_317 sky130_fd_sc_hd__decap_12
XDC_R_2_317 VGND VNB vpwr_R_317 vpwr_R_317 sky130_fd_sc_hd__decap_12
XDC_R_0_318 VGND VNB vpwr_R_318 vpwr_R_318 sky130_fd_sc_hd__decap_12
XDC_R_1_318 VGND VNB vpwr_R_318 vpwr_R_318 sky130_fd_sc_hd__decap_12
XDC_R_2_318 VGND VNB vpwr_R_318 vpwr_R_318 sky130_fd_sc_hd__decap_12
XDC_R_0_319 VGND VNB vpwr_R_319 vpwr_R_319 sky130_fd_sc_hd__decap_12
XDC_R_1_319 VGND VNB vpwr_R_319 vpwr_R_319 sky130_fd_sc_hd__decap_12
XDC_R_2_319 VGND VNB vpwr_R_319 vpwr_R_319 sky130_fd_sc_hd__decap_12
XDC_R_0_320 VGND VNB vpwr_R_320 vpwr_R_320 sky130_fd_sc_hd__decap_12
XDC_R_1_320 VGND VNB vpwr_R_320 vpwr_R_320 sky130_fd_sc_hd__decap_12
XDC_R_2_320 VGND VNB vpwr_R_320 vpwr_R_320 sky130_fd_sc_hd__decap_12
XDC_R_0_321 VGND VNB vpwr_R_321 vpwr_R_321 sky130_fd_sc_hd__decap_12
XDC_R_1_321 VGND VNB vpwr_R_321 vpwr_R_321 sky130_fd_sc_hd__decap_12
XDC_R_2_321 VGND VNB vpwr_R_321 vpwr_R_321 sky130_fd_sc_hd__decap_12
XDC_R_0_322 VGND VNB vpwr_R_322 vpwr_R_322 sky130_fd_sc_hd__decap_12
XDC_R_1_322 VGND VNB vpwr_R_322 vpwr_R_322 sky130_fd_sc_hd__decap_12
XDC_R_2_322 VGND VNB vpwr_R_322 vpwr_R_322 sky130_fd_sc_hd__decap_12
XDC_R_0_323 VGND VNB vpwr_R_323 vpwr_R_323 sky130_fd_sc_hd__decap_12
XDC_R_1_323 VGND VNB vpwr_R_323 vpwr_R_323 sky130_fd_sc_hd__decap_12
XDC_R_2_323 VGND VNB vpwr_R_323 vpwr_R_323 sky130_fd_sc_hd__decap_12
XDC_R_0_324 VGND VNB vpwr_R_324 vpwr_R_324 sky130_fd_sc_hd__decap_12
XDC_R_1_324 VGND VNB vpwr_R_324 vpwr_R_324 sky130_fd_sc_hd__decap_12
XDC_R_2_324 VGND VNB vpwr_R_324 vpwr_R_324 sky130_fd_sc_hd__decap_12
XDC_R_0_325 VGND VNB vpwr_R_325 vpwr_R_325 sky130_fd_sc_hd__decap_12
XDC_R_1_325 VGND VNB vpwr_R_325 vpwr_R_325 sky130_fd_sc_hd__decap_12
XDC_R_2_325 VGND VNB vpwr_R_325 vpwr_R_325 sky130_fd_sc_hd__decap_12
XDC_R_0_326 VGND VNB vpwr_R_326 vpwr_R_326 sky130_fd_sc_hd__decap_12
XDC_R_1_326 VGND VNB vpwr_R_326 vpwr_R_326 sky130_fd_sc_hd__decap_12
XDC_R_2_326 VGND VNB vpwr_R_326 vpwr_R_326 sky130_fd_sc_hd__decap_12
XDC_R_0_327 VGND VNB vpwr_R_327 vpwr_R_327 sky130_fd_sc_hd__decap_12
XDC_R_1_327 VGND VNB vpwr_R_327 vpwr_R_327 sky130_fd_sc_hd__decap_12
XDC_R_2_327 VGND VNB vpwr_R_327 vpwr_R_327 sky130_fd_sc_hd__decap_12
XDC_R_0_328 VGND VNB vpwr_R_328 vpwr_R_328 sky130_fd_sc_hd__decap_12
XDC_R_1_328 VGND VNB vpwr_R_328 vpwr_R_328 sky130_fd_sc_hd__decap_12
XDC_R_2_328 VGND VNB vpwr_R_328 vpwr_R_328 sky130_fd_sc_hd__decap_12
XDC_R_0_329 VGND VNB vpwr_R_329 vpwr_R_329 sky130_fd_sc_hd__decap_12
XDC_R_1_329 VGND VNB vpwr_R_329 vpwr_R_329 sky130_fd_sc_hd__decap_12
XDC_R_2_329 VGND VNB vpwr_R_329 vpwr_R_329 sky130_fd_sc_hd__decap_12
XDC_R_0_330 VGND VNB vpwr_R_330 vpwr_R_330 sky130_fd_sc_hd__decap_12
XDC_R_1_330 VGND VNB vpwr_R_330 vpwr_R_330 sky130_fd_sc_hd__decap_12
XDC_R_2_330 VGND VNB vpwr_R_330 vpwr_R_330 sky130_fd_sc_hd__decap_12
XDC_R_0_331 VGND VNB vpwr_R_331 vpwr_R_331 sky130_fd_sc_hd__decap_12
XDC_R_1_331 VGND VNB vpwr_R_331 vpwr_R_331 sky130_fd_sc_hd__decap_12
XDC_R_2_331 VGND VNB vpwr_R_331 vpwr_R_331 sky130_fd_sc_hd__decap_12
XDC_R_0_332 VGND VNB vpwr_R_332 vpwr_R_332 sky130_fd_sc_hd__decap_12
XDC_R_1_332 VGND VNB vpwr_R_332 vpwr_R_332 sky130_fd_sc_hd__decap_12
XDC_R_2_332 VGND VNB vpwr_R_332 vpwr_R_332 sky130_fd_sc_hd__decap_12
XDC_R_0_333 VGND VNB vpwr_R_333 vpwr_R_333 sky130_fd_sc_hd__decap_12
XDC_R_1_333 VGND VNB vpwr_R_333 vpwr_R_333 sky130_fd_sc_hd__decap_12
XDC_R_2_333 VGND VNB vpwr_R_333 vpwr_R_333 sky130_fd_sc_hd__decap_12
XDC_R_0_334 VGND VNB vpwr_R_334 vpwr_R_334 sky130_fd_sc_hd__decap_12
XDC_R_1_334 VGND VNB vpwr_R_334 vpwr_R_334 sky130_fd_sc_hd__decap_12
XDC_R_2_334 VGND VNB vpwr_R_334 vpwr_R_334 sky130_fd_sc_hd__decap_12
XDC_R_0_335 VGND VNB vpwr_R_335 vpwr_R_335 sky130_fd_sc_hd__decap_12
XDC_R_1_335 VGND VNB vpwr_R_335 vpwr_R_335 sky130_fd_sc_hd__decap_12
XDC_R_2_335 VGND VNB vpwr_R_335 vpwr_R_335 sky130_fd_sc_hd__decap_12
XDC_R_0_336 VGND VNB vpwr_R_336 vpwr_R_336 sky130_fd_sc_hd__decap_12
XDC_R_1_336 VGND VNB vpwr_R_336 vpwr_R_336 sky130_fd_sc_hd__decap_12
XDC_R_2_336 VGND VNB vpwr_R_336 vpwr_R_336 sky130_fd_sc_hd__decap_12
XDC_R_0_337 VGND VNB vpwr_R_337 vpwr_R_337 sky130_fd_sc_hd__decap_12
XDC_R_1_337 VGND VNB vpwr_R_337 vpwr_R_337 sky130_fd_sc_hd__decap_12
XDC_R_2_337 VGND VNB vpwr_R_337 vpwr_R_337 sky130_fd_sc_hd__decap_12
XDC_R_0_338 VGND VNB vpwr_R_338 vpwr_R_338 sky130_fd_sc_hd__decap_12
XDC_R_1_338 VGND VNB vpwr_R_338 vpwr_R_338 sky130_fd_sc_hd__decap_12
XDC_R_2_338 VGND VNB vpwr_R_338 vpwr_R_338 sky130_fd_sc_hd__decap_12
XDC_R_0_339 VGND VNB vpwr_R_339 vpwr_R_339 sky130_fd_sc_hd__decap_12
XDC_R_1_339 VGND VNB vpwr_R_339 vpwr_R_339 sky130_fd_sc_hd__decap_12
XDC_R_2_339 VGND VNB vpwr_R_339 vpwr_R_339 sky130_fd_sc_hd__decap_12
XDC_R_0_340 VGND VNB vpwr_R_340 vpwr_R_340 sky130_fd_sc_hd__decap_12
XDC_R_1_340 VGND VNB vpwr_R_340 vpwr_R_340 sky130_fd_sc_hd__decap_12
XDC_R_2_340 VGND VNB vpwr_R_340 vpwr_R_340 sky130_fd_sc_hd__decap_12
XDC_R_0_341 VGND VNB vpwr_R_341 vpwr_R_341 sky130_fd_sc_hd__decap_12
XDC_R_1_341 VGND VNB vpwr_R_341 vpwr_R_341 sky130_fd_sc_hd__decap_12
XDC_R_2_341 VGND VNB vpwr_R_341 vpwr_R_341 sky130_fd_sc_hd__decap_12
XDC_R_0_342 VGND VNB vpwr_R_342 vpwr_R_342 sky130_fd_sc_hd__decap_12
XDC_R_1_342 VGND VNB vpwr_R_342 vpwr_R_342 sky130_fd_sc_hd__decap_12
XDC_R_2_342 VGND VNB vpwr_R_342 vpwr_R_342 sky130_fd_sc_hd__decap_12
XDC_R_0_343 VGND VNB vpwr_R_343 vpwr_R_343 sky130_fd_sc_hd__decap_12
XDC_R_1_343 VGND VNB vpwr_R_343 vpwr_R_343 sky130_fd_sc_hd__decap_12
XDC_R_2_343 VGND VNB vpwr_R_343 vpwr_R_343 sky130_fd_sc_hd__decap_12
XDC_R_0_344 VGND VNB vpwr_R_344 vpwr_R_344 sky130_fd_sc_hd__decap_12
XDC_R_1_344 VGND VNB vpwr_R_344 vpwr_R_344 sky130_fd_sc_hd__decap_12
XDC_R_2_344 VGND VNB vpwr_R_344 vpwr_R_344 sky130_fd_sc_hd__decap_12
XDC_R_0_345 VGND VNB vpwr_R_345 vpwr_R_345 sky130_fd_sc_hd__decap_12
XDC_R_1_345 VGND VNB vpwr_R_345 vpwr_R_345 sky130_fd_sc_hd__decap_12
XDC_R_2_345 VGND VNB vpwr_R_345 vpwr_R_345 sky130_fd_sc_hd__decap_12
XDC_R_0_346 VGND VNB vpwr_R_346 vpwr_R_346 sky130_fd_sc_hd__decap_12
XDC_R_1_346 VGND VNB vpwr_R_346 vpwr_R_346 sky130_fd_sc_hd__decap_12
XDC_R_2_346 VGND VNB vpwr_R_346 vpwr_R_346 sky130_fd_sc_hd__decap_12
XDC_R_0_347 VGND VNB vpwr_R_347 vpwr_R_347 sky130_fd_sc_hd__decap_12
XDC_R_1_347 VGND VNB vpwr_R_347 vpwr_R_347 sky130_fd_sc_hd__decap_12
XDC_R_2_347 VGND VNB vpwr_R_347 vpwr_R_347 sky130_fd_sc_hd__decap_12
XDC_R_0_348 VGND VNB vpwr_R_348 vpwr_R_348 sky130_fd_sc_hd__decap_12
XDC_R_1_348 VGND VNB vpwr_R_348 vpwr_R_348 sky130_fd_sc_hd__decap_12
XDC_R_2_348 VGND VNB vpwr_R_348 vpwr_R_348 sky130_fd_sc_hd__decap_12
XDC_R_0_349 VGND VNB vpwr_R_349 vpwr_R_349 sky130_fd_sc_hd__decap_12
XDC_R_1_349 VGND VNB vpwr_R_349 vpwr_R_349 sky130_fd_sc_hd__decap_12
XDC_R_2_349 VGND VNB vpwr_R_349 vpwr_R_349 sky130_fd_sc_hd__decap_12
XDC_R_0_350 VGND VNB vpwr_R_350 vpwr_R_350 sky130_fd_sc_hd__decap_12
XDC_R_1_350 VGND VNB vpwr_R_350 vpwr_R_350 sky130_fd_sc_hd__decap_12
XDC_R_2_350 VGND VNB vpwr_R_350 vpwr_R_350 sky130_fd_sc_hd__decap_12
XDC_R_0_351 VGND VNB vpwr_R_351 vpwr_R_351 sky130_fd_sc_hd__decap_12
XDC_R_1_351 VGND VNB vpwr_R_351 vpwr_R_351 sky130_fd_sc_hd__decap_12
XDC_R_2_351 VGND VNB vpwr_R_351 vpwr_R_351 sky130_fd_sc_hd__decap_12
XDC_R_0_352 VGND VNB vpwr_R_352 vpwr_R_352 sky130_fd_sc_hd__decap_12
XDC_R_1_352 VGND VNB vpwr_R_352 vpwr_R_352 sky130_fd_sc_hd__decap_12
XDC_R_2_352 VGND VNB vpwr_R_352 vpwr_R_352 sky130_fd_sc_hd__decap_12
XDC_R_0_353 VGND VNB vpwr_R_353 vpwr_R_353 sky130_fd_sc_hd__decap_12
XDC_R_1_353 VGND VNB vpwr_R_353 vpwr_R_353 sky130_fd_sc_hd__decap_12
XDC_R_2_353 VGND VNB vpwr_R_353 vpwr_R_353 sky130_fd_sc_hd__decap_12
XDC_R_0_354 VGND VNB vpwr_R_354 vpwr_R_354 sky130_fd_sc_hd__decap_12
XDC_R_1_354 VGND VNB vpwr_R_354 vpwr_R_354 sky130_fd_sc_hd__decap_12
XDC_R_2_354 VGND VNB vpwr_R_354 vpwr_R_354 sky130_fd_sc_hd__decap_12
XDC_R_0_355 VGND VNB vpwr_R_355 vpwr_R_355 sky130_fd_sc_hd__decap_12
XDC_R_1_355 VGND VNB vpwr_R_355 vpwr_R_355 sky130_fd_sc_hd__decap_12
XDC_R_2_355 VGND VNB vpwr_R_355 vpwr_R_355 sky130_fd_sc_hd__decap_12
XDC_R_0_356 VGND VNB vpwr_R_356 vpwr_R_356 sky130_fd_sc_hd__decap_12
XDC_R_1_356 VGND VNB vpwr_R_356 vpwr_R_356 sky130_fd_sc_hd__decap_12
XDC_R_2_356 VGND VNB vpwr_R_356 vpwr_R_356 sky130_fd_sc_hd__decap_12
XDC_R_0_357 VGND VNB vpwr_R_357 vpwr_R_357 sky130_fd_sc_hd__decap_12
XDC_R_1_357 VGND VNB vpwr_R_357 vpwr_R_357 sky130_fd_sc_hd__decap_12
XDC_R_2_357 VGND VNB vpwr_R_357 vpwr_R_357 sky130_fd_sc_hd__decap_12
XDC_R_0_358 VGND VNB vpwr_R_358 vpwr_R_358 sky130_fd_sc_hd__decap_12
XDC_R_1_358 VGND VNB vpwr_R_358 vpwr_R_358 sky130_fd_sc_hd__decap_12
XDC_R_2_358 VGND VNB vpwr_R_358 vpwr_R_358 sky130_fd_sc_hd__decap_12
XDC_R_0_359 VGND VNB vpwr_R_359 vpwr_R_359 sky130_fd_sc_hd__decap_12
XDC_R_1_359 VGND VNB vpwr_R_359 vpwr_R_359 sky130_fd_sc_hd__decap_12
XDC_R_2_359 VGND VNB vpwr_R_359 vpwr_R_359 sky130_fd_sc_hd__decap_12
XDC_R_0_360 VGND VNB vpwr_R_360 vpwr_R_360 sky130_fd_sc_hd__decap_12
XDC_R_1_360 VGND VNB vpwr_R_360 vpwr_R_360 sky130_fd_sc_hd__decap_12
XDC_R_2_360 VGND VNB vpwr_R_360 vpwr_R_360 sky130_fd_sc_hd__decap_12
XDC_R_0_361 VGND VNB vpwr_R_361 vpwr_R_361 sky130_fd_sc_hd__decap_12
XDC_R_1_361 VGND VNB vpwr_R_361 vpwr_R_361 sky130_fd_sc_hd__decap_12
XDC_R_2_361 VGND VNB vpwr_R_361 vpwr_R_361 sky130_fd_sc_hd__decap_12
XDC_R_0_362 VGND VNB vpwr_R_362 vpwr_R_362 sky130_fd_sc_hd__decap_12
XDC_R_1_362 VGND VNB vpwr_R_362 vpwr_R_362 sky130_fd_sc_hd__decap_12
XDC_R_2_362 VGND VNB vpwr_R_362 vpwr_R_362 sky130_fd_sc_hd__decap_12
XDC_R_0_363 VGND VNB vpwr_R_363 vpwr_R_363 sky130_fd_sc_hd__decap_12
XDC_R_1_363 VGND VNB vpwr_R_363 vpwr_R_363 sky130_fd_sc_hd__decap_12
XDC_R_2_363 VGND VNB vpwr_R_363 vpwr_R_363 sky130_fd_sc_hd__decap_12
XDC_R_0_364 VGND VNB vpwr_R_364 vpwr_R_364 sky130_fd_sc_hd__decap_12
XDC_R_1_364 VGND VNB vpwr_R_364 vpwr_R_364 sky130_fd_sc_hd__decap_12
XDC_R_2_364 VGND VNB vpwr_R_364 vpwr_R_364 sky130_fd_sc_hd__decap_12
XDC_R_0_365 VGND VNB vpwr_R_365 vpwr_R_365 sky130_fd_sc_hd__decap_12
XDC_R_1_365 VGND VNB vpwr_R_365 vpwr_R_365 sky130_fd_sc_hd__decap_12
XDC_R_2_365 VGND VNB vpwr_R_365 vpwr_R_365 sky130_fd_sc_hd__decap_12
XDC_R_0_366 VGND VNB vpwr_R_366 vpwr_R_366 sky130_fd_sc_hd__decap_12
XDC_R_1_366 VGND VNB vpwr_R_366 vpwr_R_366 sky130_fd_sc_hd__decap_12
XDC_R_2_366 VGND VNB vpwr_R_366 vpwr_R_366 sky130_fd_sc_hd__decap_12
XDC_R_0_367 VGND VNB vpwr_R_367 vpwr_R_367 sky130_fd_sc_hd__decap_12
XDC_R_1_367 VGND VNB vpwr_R_367 vpwr_R_367 sky130_fd_sc_hd__decap_12
XDC_R_2_367 VGND VNB vpwr_R_367 vpwr_R_367 sky130_fd_sc_hd__decap_12
XDC_R_0_368 VGND VNB vpwr_R_368 vpwr_R_368 sky130_fd_sc_hd__decap_12
XDC_R_1_368 VGND VNB vpwr_R_368 vpwr_R_368 sky130_fd_sc_hd__decap_12
XDC_R_2_368 VGND VNB vpwr_R_368 vpwr_R_368 sky130_fd_sc_hd__decap_12
XDC_R_0_369 VGND VNB vpwr_R_369 vpwr_R_369 sky130_fd_sc_hd__decap_12
XDC_R_1_369 VGND VNB vpwr_R_369 vpwr_R_369 sky130_fd_sc_hd__decap_12
XDC_R_2_369 VGND VNB vpwr_R_369 vpwr_R_369 sky130_fd_sc_hd__decap_12
XDC_R_0_370 VGND VNB vpwr_R_370 vpwr_R_370 sky130_fd_sc_hd__decap_12
XDC_R_1_370 VGND VNB vpwr_R_370 vpwr_R_370 sky130_fd_sc_hd__decap_12
XDC_R_2_370 VGND VNB vpwr_R_370 vpwr_R_370 sky130_fd_sc_hd__decap_12
XDC_R_0_371 VGND VNB vpwr_R_371 vpwr_R_371 sky130_fd_sc_hd__decap_12
XDC_R_1_371 VGND VNB vpwr_R_371 vpwr_R_371 sky130_fd_sc_hd__decap_12
XDC_R_2_371 VGND VNB vpwr_R_371 vpwr_R_371 sky130_fd_sc_hd__decap_12
XDC_R_0_372 VGND VNB vpwr_R_372 vpwr_R_372 sky130_fd_sc_hd__decap_12
XDC_R_1_372 VGND VNB vpwr_R_372 vpwr_R_372 sky130_fd_sc_hd__decap_12
XDC_R_2_372 VGND VNB vpwr_R_372 vpwr_R_372 sky130_fd_sc_hd__decap_12
XDC_R_0_373 VGND VNB vpwr_R_373 vpwr_R_373 sky130_fd_sc_hd__decap_12
XDC_R_1_373 VGND VNB vpwr_R_373 vpwr_R_373 sky130_fd_sc_hd__decap_12
XDC_R_2_373 VGND VNB vpwr_R_373 vpwr_R_373 sky130_fd_sc_hd__decap_12
XDC_R_0_374 VGND VNB vpwr_R_374 vpwr_R_374 sky130_fd_sc_hd__decap_12
XDC_R_1_374 VGND VNB vpwr_R_374 vpwr_R_374 sky130_fd_sc_hd__decap_12
XDC_R_2_374 VGND VNB vpwr_R_374 vpwr_R_374 sky130_fd_sc_hd__decap_12
XDC_R_0_375 VGND VNB vpwr_R_375 vpwr_R_375 sky130_fd_sc_hd__decap_12
XDC_R_1_375 VGND VNB vpwr_R_375 vpwr_R_375 sky130_fd_sc_hd__decap_12
XDC_R_2_375 VGND VNB vpwr_R_375 vpwr_R_375 sky130_fd_sc_hd__decap_12
XDC_R_0_376 VGND VNB vpwr_R_376 vpwr_R_376 sky130_fd_sc_hd__decap_12
XDC_R_1_376 VGND VNB vpwr_R_376 vpwr_R_376 sky130_fd_sc_hd__decap_12
XDC_R_2_376 VGND VNB vpwr_R_376 vpwr_R_376 sky130_fd_sc_hd__decap_12
XDC_R_0_377 VGND VNB vpwr_R_377 vpwr_R_377 sky130_fd_sc_hd__decap_12
XDC_R_1_377 VGND VNB vpwr_R_377 vpwr_R_377 sky130_fd_sc_hd__decap_12
XDC_R_2_377 VGND VNB vpwr_R_377 vpwr_R_377 sky130_fd_sc_hd__decap_12
XDC_R_0_378 VGND VNB vpwr_R_378 vpwr_R_378 sky130_fd_sc_hd__decap_12
XDC_R_1_378 VGND VNB vpwr_R_378 vpwr_R_378 sky130_fd_sc_hd__decap_12
XDC_R_2_378 VGND VNB vpwr_R_378 vpwr_R_378 sky130_fd_sc_hd__decap_12
XDC_R_0_379 VGND VNB vpwr_R_379 vpwr_R_379 sky130_fd_sc_hd__decap_12
XDC_R_1_379 VGND VNB vpwr_R_379 vpwr_R_379 sky130_fd_sc_hd__decap_12
XDC_R_2_379 VGND VNB vpwr_R_379 vpwr_R_379 sky130_fd_sc_hd__decap_12
XDC_R_0_380 VGND VNB vpwr_R_380 vpwr_R_380 sky130_fd_sc_hd__decap_12
XDC_R_1_380 VGND VNB vpwr_R_380 vpwr_R_380 sky130_fd_sc_hd__decap_12
XDC_R_2_380 VGND VNB vpwr_R_380 vpwr_R_380 sky130_fd_sc_hd__decap_12
XDC_R_0_381 VGND VNB vpwr_R_381 vpwr_R_381 sky130_fd_sc_hd__decap_12
XDC_R_1_381 VGND VNB vpwr_R_381 vpwr_R_381 sky130_fd_sc_hd__decap_12
XDC_R_2_381 VGND VNB vpwr_R_381 vpwr_R_381 sky130_fd_sc_hd__decap_12
XDC_R_0_382 VGND VNB vpwr_R_382 vpwr_R_382 sky130_fd_sc_hd__decap_12
XDC_R_1_382 VGND VNB vpwr_R_382 vpwr_R_382 sky130_fd_sc_hd__decap_12
XDC_R_2_382 VGND VNB vpwr_R_382 vpwr_R_382 sky130_fd_sc_hd__decap_12
XDC_R_0_383 VGND VNB vpwr_R_383 vpwr_R_383 sky130_fd_sc_hd__decap_12
XDC_R_1_383 VGND VNB vpwr_R_383 vpwr_R_383 sky130_fd_sc_hd__decap_12
XDC_R_2_383 VGND VNB vpwr_R_383 vpwr_R_383 sky130_fd_sc_hd__decap_12
XDC_R_0_384 VGND VNB vpwr_R_384 vpwr_R_384 sky130_fd_sc_hd__decap_12
XDC_R_1_384 VGND VNB vpwr_R_384 vpwr_R_384 sky130_fd_sc_hd__decap_12
XDC_R_2_384 VGND VNB vpwr_R_384 vpwr_R_384 sky130_fd_sc_hd__decap_12
XDC_R_0_385 VGND VNB vpwr_R_385 vpwr_R_385 sky130_fd_sc_hd__decap_12
XDC_R_1_385 VGND VNB vpwr_R_385 vpwr_R_385 sky130_fd_sc_hd__decap_12
XDC_R_2_385 VGND VNB vpwr_R_385 vpwr_R_385 sky130_fd_sc_hd__decap_12
XDC_R_0_386 VGND VNB vpwr_R_386 vpwr_R_386 sky130_fd_sc_hd__decap_12
XDC_R_1_386 VGND VNB vpwr_R_386 vpwr_R_386 sky130_fd_sc_hd__decap_12
XDC_R_2_386 VGND VNB vpwr_R_386 vpwr_R_386 sky130_fd_sc_hd__decap_12
XDC_R_0_387 VGND VNB vpwr_R_387 vpwr_R_387 sky130_fd_sc_hd__decap_12
XDC_R_1_387 VGND VNB vpwr_R_387 vpwr_R_387 sky130_fd_sc_hd__decap_12
XDC_R_2_387 VGND VNB vpwr_R_387 vpwr_R_387 sky130_fd_sc_hd__decap_12
XDC_R_0_388 VGND VNB vpwr_R_388 vpwr_R_388 sky130_fd_sc_hd__decap_12
XDC_R_1_388 VGND VNB vpwr_R_388 vpwr_R_388 sky130_fd_sc_hd__decap_12
XDC_R_2_388 VGND VNB vpwr_R_388 vpwr_R_388 sky130_fd_sc_hd__decap_12
XDC_R_0_389 VGND VNB vpwr_R_389 vpwr_R_389 sky130_fd_sc_hd__decap_12
XDC_R_1_389 VGND VNB vpwr_R_389 vpwr_R_389 sky130_fd_sc_hd__decap_12
XDC_R_2_389 VGND VNB vpwr_R_389 vpwr_R_389 sky130_fd_sc_hd__decap_12
XDC_R_0_390 VGND VNB vpwr_R_390 vpwr_R_390 sky130_fd_sc_hd__decap_12
XDC_R_1_390 VGND VNB vpwr_R_390 vpwr_R_390 sky130_fd_sc_hd__decap_12
XDC_R_2_390 VGND VNB vpwr_R_390 vpwr_R_390 sky130_fd_sc_hd__decap_12
XDC_R_0_391 VGND VNB vpwr_R_391 vpwr_R_391 sky130_fd_sc_hd__decap_12
XDC_R_1_391 VGND VNB vpwr_R_391 vpwr_R_391 sky130_fd_sc_hd__decap_12
XDC_R_2_391 VGND VNB vpwr_R_391 vpwr_R_391 sky130_fd_sc_hd__decap_12
XDC_R_0_392 VGND VNB vpwr_R_392 vpwr_R_392 sky130_fd_sc_hd__decap_12
XDC_R_1_392 VGND VNB vpwr_R_392 vpwr_R_392 sky130_fd_sc_hd__decap_12
XDC_R_2_392 VGND VNB vpwr_R_392 vpwr_R_392 sky130_fd_sc_hd__decap_12
XDC_R_0_393 VGND VNB vpwr_R_393 vpwr_R_393 sky130_fd_sc_hd__decap_12
XDC_R_1_393 VGND VNB vpwr_R_393 vpwr_R_393 sky130_fd_sc_hd__decap_12
XDC_R_2_393 VGND VNB vpwr_R_393 vpwr_R_393 sky130_fd_sc_hd__decap_12
XDC_R_0_394 VGND VNB vpwr_R_394 vpwr_R_394 sky130_fd_sc_hd__decap_12
XDC_R_1_394 VGND VNB vpwr_R_394 vpwr_R_394 sky130_fd_sc_hd__decap_12
XDC_R_2_394 VGND VNB vpwr_R_394 vpwr_R_394 sky130_fd_sc_hd__decap_12
XDC_R_0_395 VGND VNB vpwr_R_395 vpwr_R_395 sky130_fd_sc_hd__decap_12
XDC_R_1_395 VGND VNB vpwr_R_395 vpwr_R_395 sky130_fd_sc_hd__decap_12
XDC_R_2_395 VGND VNB vpwr_R_395 vpwr_R_395 sky130_fd_sc_hd__decap_12
XDC_R_0_396 VGND VNB vpwr_R_396 vpwr_R_396 sky130_fd_sc_hd__decap_12
XDC_R_1_396 VGND VNB vpwr_R_396 vpwr_R_396 sky130_fd_sc_hd__decap_12
XDC_R_2_396 VGND VNB vpwr_R_396 vpwr_R_396 sky130_fd_sc_hd__decap_12
XDC_R_0_397 VGND VNB vpwr_R_397 vpwr_R_397 sky130_fd_sc_hd__decap_12
XDC_R_1_397 VGND VNB vpwr_R_397 vpwr_R_397 sky130_fd_sc_hd__decap_12
XDC_R_2_397 VGND VNB vpwr_R_397 vpwr_R_397 sky130_fd_sc_hd__decap_12
XDC_R_0_398 VGND VNB vpwr_R_398 vpwr_R_398 sky130_fd_sc_hd__decap_12
XDC_R_1_398 VGND VNB vpwr_R_398 vpwr_R_398 sky130_fd_sc_hd__decap_12
XDC_R_2_398 VGND VNB vpwr_R_398 vpwr_R_398 sky130_fd_sc_hd__decap_12
XDC_R_0_399 VGND VNB vpwr_R_399 vpwr_R_399 sky130_fd_sc_hd__decap_12
XDC_R_1_399 VGND VNB vpwr_R_399 vpwr_R_399 sky130_fd_sc_hd__decap_12
XDC_R_2_399 VGND VNB vpwr_R_399 vpwr_R_399 sky130_fd_sc_hd__decap_12
XDC_R_0_400 VGND VNB vpwr_R_400 vpwr_R_400 sky130_fd_sc_hd__decap_12
XDC_R_1_400 VGND VNB vpwr_R_400 vpwr_R_400 sky130_fd_sc_hd__decap_12
XDC_R_2_400 VGND VNB vpwr_R_400 vpwr_R_400 sky130_fd_sc_hd__decap_12
XDC_R_0_401 VGND VNB vpwr_R_401 vpwr_R_401 sky130_fd_sc_hd__decap_12
XDC_R_1_401 VGND VNB vpwr_R_401 vpwr_R_401 sky130_fd_sc_hd__decap_12
XDC_R_2_401 VGND VNB vpwr_R_401 vpwr_R_401 sky130_fd_sc_hd__decap_12
XDC_R_0_402 VGND VNB vpwr_R_402 vpwr_R_402 sky130_fd_sc_hd__decap_12
XDC_R_1_402 VGND VNB vpwr_R_402 vpwr_R_402 sky130_fd_sc_hd__decap_12
XDC_R_2_402 VGND VNB vpwr_R_402 vpwr_R_402 sky130_fd_sc_hd__decap_12
XDC_R_0_403 VGND VNB vpwr_R_403 vpwr_R_403 sky130_fd_sc_hd__decap_12
XDC_R_1_403 VGND VNB vpwr_R_403 vpwr_R_403 sky130_fd_sc_hd__decap_12
XDC_R_2_403 VGND VNB vpwr_R_403 vpwr_R_403 sky130_fd_sc_hd__decap_12
XDC_R_0_404 VGND VNB vpwr_R_404 vpwr_R_404 sky130_fd_sc_hd__decap_12
XDC_R_1_404 VGND VNB vpwr_R_404 vpwr_R_404 sky130_fd_sc_hd__decap_12
XDC_R_2_404 VGND VNB vpwr_R_404 vpwr_R_404 sky130_fd_sc_hd__decap_12
XDC_R_0_405 VGND VNB vpwr_R_405 vpwr_R_405 sky130_fd_sc_hd__decap_12
XDC_R_1_405 VGND VNB vpwr_R_405 vpwr_R_405 sky130_fd_sc_hd__decap_12
XDC_R_2_405 VGND VNB vpwr_R_405 vpwr_R_405 sky130_fd_sc_hd__decap_12
XDC_R_0_406 VGND VNB vpwr_R_406 vpwr_R_406 sky130_fd_sc_hd__decap_12
XDC_R_1_406 VGND VNB vpwr_R_406 vpwr_R_406 sky130_fd_sc_hd__decap_12
XDC_R_2_406 VGND VNB vpwr_R_406 vpwr_R_406 sky130_fd_sc_hd__decap_12
XDC_R_0_407 VGND VNB vpwr_R_407 vpwr_R_407 sky130_fd_sc_hd__decap_12
XDC_R_1_407 VGND VNB vpwr_R_407 vpwr_R_407 sky130_fd_sc_hd__decap_12
XDC_R_2_407 VGND VNB vpwr_R_407 vpwr_R_407 sky130_fd_sc_hd__decap_12
XDC_R_0_408 VGND VNB vpwr_R_408 vpwr_R_408 sky130_fd_sc_hd__decap_12
XDC_R_1_408 VGND VNB vpwr_R_408 vpwr_R_408 sky130_fd_sc_hd__decap_12
XDC_R_2_408 VGND VNB vpwr_R_408 vpwr_R_408 sky130_fd_sc_hd__decap_12
XDC_R_0_409 VGND VNB vpwr_R_409 vpwr_R_409 sky130_fd_sc_hd__decap_12
XDC_R_1_409 VGND VNB vpwr_R_409 vpwr_R_409 sky130_fd_sc_hd__decap_12
XDC_R_2_409 VGND VNB vpwr_R_409 vpwr_R_409 sky130_fd_sc_hd__decap_12
XDC_R_0_410 VGND VNB vpwr_R_410 vpwr_R_410 sky130_fd_sc_hd__decap_12
XDC_R_1_410 VGND VNB vpwr_R_410 vpwr_R_410 sky130_fd_sc_hd__decap_12
XDC_R_2_410 VGND VNB vpwr_R_410 vpwr_R_410 sky130_fd_sc_hd__decap_12
XDC_R_0_411 VGND VNB vpwr_R_411 vpwr_R_411 sky130_fd_sc_hd__decap_12
XDC_R_1_411 VGND VNB vpwr_R_411 vpwr_R_411 sky130_fd_sc_hd__decap_12
XDC_R_2_411 VGND VNB vpwr_R_411 vpwr_R_411 sky130_fd_sc_hd__decap_12
XDC_R_0_412 VGND VNB vpwr_R_412 vpwr_R_412 sky130_fd_sc_hd__decap_12
XDC_R_1_412 VGND VNB vpwr_R_412 vpwr_R_412 sky130_fd_sc_hd__decap_12
XDC_R_2_412 VGND VNB vpwr_R_412 vpwr_R_412 sky130_fd_sc_hd__decap_12
XDC_R_0_413 VGND VNB vpwr_R_413 vpwr_R_413 sky130_fd_sc_hd__decap_12
XDC_R_1_413 VGND VNB vpwr_R_413 vpwr_R_413 sky130_fd_sc_hd__decap_12
XDC_R_2_413 VGND VNB vpwr_R_413 vpwr_R_413 sky130_fd_sc_hd__decap_12
XDC_R_0_414 VGND VNB vpwr_R_414 vpwr_R_414 sky130_fd_sc_hd__decap_12
XDC_R_1_414 VGND VNB vpwr_R_414 vpwr_R_414 sky130_fd_sc_hd__decap_12
XDC_R_2_414 VGND VNB vpwr_R_414 vpwr_R_414 sky130_fd_sc_hd__decap_12
XDC_R_0_415 VGND VNB vpwr_R_415 vpwr_R_415 sky130_fd_sc_hd__decap_12
XDC_R_1_415 VGND VNB vpwr_R_415 vpwr_R_415 sky130_fd_sc_hd__decap_12
XDC_R_2_415 VGND VNB vpwr_R_415 vpwr_R_415 sky130_fd_sc_hd__decap_12
XDC_R_0_416 VGND VNB vpwr_R_416 vpwr_R_416 sky130_fd_sc_hd__decap_12
XDC_R_1_416 VGND VNB vpwr_R_416 vpwr_R_416 sky130_fd_sc_hd__decap_12
XDC_R_2_416 VGND VNB vpwr_R_416 vpwr_R_416 sky130_fd_sc_hd__decap_12
XDC_R_0_417 VGND VNB vpwr_R_417 vpwr_R_417 sky130_fd_sc_hd__decap_12
XDC_R_1_417 VGND VNB vpwr_R_417 vpwr_R_417 sky130_fd_sc_hd__decap_12
XDC_R_2_417 VGND VNB vpwr_R_417 vpwr_R_417 sky130_fd_sc_hd__decap_12
XDC_R_0_418 VGND VNB vpwr_R_418 vpwr_R_418 sky130_fd_sc_hd__decap_12
XDC_R_1_418 VGND VNB vpwr_R_418 vpwr_R_418 sky130_fd_sc_hd__decap_12
XDC_R_2_418 VGND VNB vpwr_R_418 vpwr_R_418 sky130_fd_sc_hd__decap_12
XDC_R_0_419 VGND VNB vpwr_R_419 vpwr_R_419 sky130_fd_sc_hd__decap_12
XDC_R_1_419 VGND VNB vpwr_R_419 vpwr_R_419 sky130_fd_sc_hd__decap_12
XDC_R_2_419 VGND VNB vpwr_R_419 vpwr_R_419 sky130_fd_sc_hd__decap_12
XDC_R_0_420 VGND VNB vpwr_R_420 vpwr_R_420 sky130_fd_sc_hd__decap_12
XDC_R_1_420 VGND VNB vpwr_R_420 vpwr_R_420 sky130_fd_sc_hd__decap_12
XDC_R_2_420 VGND VNB vpwr_R_420 vpwr_R_420 sky130_fd_sc_hd__decap_12
XDC_R_0_421 VGND VNB vpwr_R_421 vpwr_R_421 sky130_fd_sc_hd__decap_12
XDC_R_1_421 VGND VNB vpwr_R_421 vpwr_R_421 sky130_fd_sc_hd__decap_12
XDC_R_2_421 VGND VNB vpwr_R_421 vpwr_R_421 sky130_fd_sc_hd__decap_12
XDC_R_0_422 VGND VNB vpwr_R_422 vpwr_R_422 sky130_fd_sc_hd__decap_12
XDC_R_1_422 VGND VNB vpwr_R_422 vpwr_R_422 sky130_fd_sc_hd__decap_12
XDC_R_2_422 VGND VNB vpwr_R_422 vpwr_R_422 sky130_fd_sc_hd__decap_12
XDC_R_0_423 VGND VNB vpwr_R_423 vpwr_R_423 sky130_fd_sc_hd__decap_12
XDC_R_1_423 VGND VNB vpwr_R_423 vpwr_R_423 sky130_fd_sc_hd__decap_12
XDC_R_2_423 VGND VNB vpwr_R_423 vpwr_R_423 sky130_fd_sc_hd__decap_12
XDC_R_0_424 VGND VNB vpwr_R_424 vpwr_R_424 sky130_fd_sc_hd__decap_12
XDC_R_1_424 VGND VNB vpwr_R_424 vpwr_R_424 sky130_fd_sc_hd__decap_12
XDC_R_2_424 VGND VNB vpwr_R_424 vpwr_R_424 sky130_fd_sc_hd__decap_12
XDC_R_0_425 VGND VNB vpwr_R_425 vpwr_R_425 sky130_fd_sc_hd__decap_12
XDC_R_1_425 VGND VNB vpwr_R_425 vpwr_R_425 sky130_fd_sc_hd__decap_12
XDC_R_2_425 VGND VNB vpwr_R_425 vpwr_R_425 sky130_fd_sc_hd__decap_12
XDC_R_0_426 VGND VNB vpwr_R_426 vpwr_R_426 sky130_fd_sc_hd__decap_12
XDC_R_1_426 VGND VNB vpwr_R_426 vpwr_R_426 sky130_fd_sc_hd__decap_12
XDC_R_2_426 VGND VNB vpwr_R_426 vpwr_R_426 sky130_fd_sc_hd__decap_12
XDC_R_0_427 VGND VNB vpwr_R_427 vpwr_R_427 sky130_fd_sc_hd__decap_12
XDC_R_1_427 VGND VNB vpwr_R_427 vpwr_R_427 sky130_fd_sc_hd__decap_12
XDC_R_2_427 VGND VNB vpwr_R_427 vpwr_R_427 sky130_fd_sc_hd__decap_12
XDC_R_0_428 VGND VNB vpwr_R_428 vpwr_R_428 sky130_fd_sc_hd__decap_12
XDC_R_1_428 VGND VNB vpwr_R_428 vpwr_R_428 sky130_fd_sc_hd__decap_12
XDC_R_2_428 VGND VNB vpwr_R_428 vpwr_R_428 sky130_fd_sc_hd__decap_12
XDC_R_0_429 VGND VNB vpwr_R_429 vpwr_R_429 sky130_fd_sc_hd__decap_12
XDC_R_1_429 VGND VNB vpwr_R_429 vpwr_R_429 sky130_fd_sc_hd__decap_12
XDC_R_2_429 VGND VNB vpwr_R_429 vpwr_R_429 sky130_fd_sc_hd__decap_12
XDC_R_0_430 VGND VNB vpwr_R_430 vpwr_R_430 sky130_fd_sc_hd__decap_12
XDC_R_1_430 VGND VNB vpwr_R_430 vpwr_R_430 sky130_fd_sc_hd__decap_12
XDC_R_2_430 VGND VNB vpwr_R_430 vpwr_R_430 sky130_fd_sc_hd__decap_12
XDC_R_0_431 VGND VNB vpwr_R_431 vpwr_R_431 sky130_fd_sc_hd__decap_12
XDC_R_1_431 VGND VNB vpwr_R_431 vpwr_R_431 sky130_fd_sc_hd__decap_12
XDC_R_2_431 VGND VNB vpwr_R_431 vpwr_R_431 sky130_fd_sc_hd__decap_12
XDC_R_0_432 VGND VNB vpwr_R_432 vpwr_R_432 sky130_fd_sc_hd__decap_12
XDC_R_1_432 VGND VNB vpwr_R_432 vpwr_R_432 sky130_fd_sc_hd__decap_12
XDC_R_2_432 VGND VNB vpwr_R_432 vpwr_R_432 sky130_fd_sc_hd__decap_12
XDC_R_0_433 VGND VNB vpwr_R_433 vpwr_R_433 sky130_fd_sc_hd__decap_12
XDC_R_1_433 VGND VNB vpwr_R_433 vpwr_R_433 sky130_fd_sc_hd__decap_12
XDC_R_2_433 VGND VNB vpwr_R_433 vpwr_R_433 sky130_fd_sc_hd__decap_12
XDC_R_0_434 VGND VNB vpwr_R_434 vpwr_R_434 sky130_fd_sc_hd__decap_12
XDC_R_1_434 VGND VNB vpwr_R_434 vpwr_R_434 sky130_fd_sc_hd__decap_12
XDC_R_2_434 VGND VNB vpwr_R_434 vpwr_R_434 sky130_fd_sc_hd__decap_12
XDC_R_0_435 VGND VNB vpwr_R_435 vpwr_R_435 sky130_fd_sc_hd__decap_12
XDC_R_1_435 VGND VNB vpwr_R_435 vpwr_R_435 sky130_fd_sc_hd__decap_12
XDC_R_2_435 VGND VNB vpwr_R_435 vpwr_R_435 sky130_fd_sc_hd__decap_12
XDC_R_0_436 VGND VNB vpwr_R_436 vpwr_R_436 sky130_fd_sc_hd__decap_12
XDC_R_1_436 VGND VNB vpwr_R_436 vpwr_R_436 sky130_fd_sc_hd__decap_12
XDC_R_2_436 VGND VNB vpwr_R_436 vpwr_R_436 sky130_fd_sc_hd__decap_12
XDC_R_0_437 VGND VNB vpwr_R_437 vpwr_R_437 sky130_fd_sc_hd__decap_12
XDC_R_1_437 VGND VNB vpwr_R_437 vpwr_R_437 sky130_fd_sc_hd__decap_12
XDC_R_2_437 VGND VNB vpwr_R_437 vpwr_R_437 sky130_fd_sc_hd__decap_12
XDC_R_0_438 VGND VNB vpwr_R_438 vpwr_R_438 sky130_fd_sc_hd__decap_12
XDC_R_1_438 VGND VNB vpwr_R_438 vpwr_R_438 sky130_fd_sc_hd__decap_12
XDC_R_2_438 VGND VNB vpwr_R_438 vpwr_R_438 sky130_fd_sc_hd__decap_12
XDC_R_0_439 VGND VNB vpwr_R_439 vpwr_R_439 sky130_fd_sc_hd__decap_12
XDC_R_1_439 VGND VNB vpwr_R_439 vpwr_R_439 sky130_fd_sc_hd__decap_12
XDC_R_2_439 VGND VNB vpwr_R_439 vpwr_R_439 sky130_fd_sc_hd__decap_12
XDC_R_0_440 VGND VNB vpwr_R_440 vpwr_R_440 sky130_fd_sc_hd__decap_12
XDC_R_1_440 VGND VNB vpwr_R_440 vpwr_R_440 sky130_fd_sc_hd__decap_12
XDC_R_2_440 VGND VNB vpwr_R_440 vpwr_R_440 sky130_fd_sc_hd__decap_12
XDC_R_0_441 VGND VNB vpwr_R_441 vpwr_R_441 sky130_fd_sc_hd__decap_12
XDC_R_1_441 VGND VNB vpwr_R_441 vpwr_R_441 sky130_fd_sc_hd__decap_12
XDC_R_2_441 VGND VNB vpwr_R_441 vpwr_R_441 sky130_fd_sc_hd__decap_12
XDC_R_0_442 VGND VNB vpwr_R_442 vpwr_R_442 sky130_fd_sc_hd__decap_12
XDC_R_1_442 VGND VNB vpwr_R_442 vpwr_R_442 sky130_fd_sc_hd__decap_12
XDC_R_2_442 VGND VNB vpwr_R_442 vpwr_R_442 sky130_fd_sc_hd__decap_12
XDC_R_0_443 VGND VNB vpwr_R_443 vpwr_R_443 sky130_fd_sc_hd__decap_12
XDC_R_1_443 VGND VNB vpwr_R_443 vpwr_R_443 sky130_fd_sc_hd__decap_12
XDC_R_2_443 VGND VNB vpwr_R_443 vpwr_R_443 sky130_fd_sc_hd__decap_12
XDC_R_0_444 VGND VNB vpwr_R_444 vpwr_R_444 sky130_fd_sc_hd__decap_12
XDC_R_1_444 VGND VNB vpwr_R_444 vpwr_R_444 sky130_fd_sc_hd__decap_12
XDC_R_2_444 VGND VNB vpwr_R_444 vpwr_R_444 sky130_fd_sc_hd__decap_12
XDC_R_0_445 VGND VNB vpwr_R_445 vpwr_R_445 sky130_fd_sc_hd__decap_12
XDC_R_1_445 VGND VNB vpwr_R_445 vpwr_R_445 sky130_fd_sc_hd__decap_12
XDC_R_2_445 VGND VNB vpwr_R_445 vpwr_R_445 sky130_fd_sc_hd__decap_12
XDC_R_0_446 VGND VNB vpwr_R_446 vpwr_R_446 sky130_fd_sc_hd__decap_12
XDC_R_1_446 VGND VNB vpwr_R_446 vpwr_R_446 sky130_fd_sc_hd__decap_12
XDC_R_2_446 VGND VNB vpwr_R_446 vpwr_R_446 sky130_fd_sc_hd__decap_12
XDC_R_0_447 VGND VNB vpwr_R_447 vpwr_R_447 sky130_fd_sc_hd__decap_12
XDC_R_1_447 VGND VNB vpwr_R_447 vpwr_R_447 sky130_fd_sc_hd__decap_12
XDC_R_2_447 VGND VNB vpwr_R_447 vpwr_R_447 sky130_fd_sc_hd__decap_12
XDC_R_0_448 VGND VNB vpwr_R_448 vpwr_R_448 sky130_fd_sc_hd__decap_12
XDC_R_1_448 VGND VNB vpwr_R_448 vpwr_R_448 sky130_fd_sc_hd__decap_12
XDC_R_2_448 VGND VNB vpwr_R_448 vpwr_R_448 sky130_fd_sc_hd__decap_12
XDC_R_0_449 VGND VNB vpwr_R_449 vpwr_R_449 sky130_fd_sc_hd__decap_12
XDC_R_1_449 VGND VNB vpwr_R_449 vpwr_R_449 sky130_fd_sc_hd__decap_12
XDC_R_2_449 VGND VNB vpwr_R_449 vpwr_R_449 sky130_fd_sc_hd__decap_12
XDC_R_0_450 VGND VNB vpwr_R_450 vpwr_R_450 sky130_fd_sc_hd__decap_12
XDC_R_1_450 VGND VNB vpwr_R_450 vpwr_R_450 sky130_fd_sc_hd__decap_12
XDC_R_2_450 VGND VNB vpwr_R_450 vpwr_R_450 sky130_fd_sc_hd__decap_12
XDC_R_0_451 VGND VNB vpwr_R_451 vpwr_R_451 sky130_fd_sc_hd__decap_12
XDC_R_1_451 VGND VNB vpwr_R_451 vpwr_R_451 sky130_fd_sc_hd__decap_12
XDC_R_2_451 VGND VNB vpwr_R_451 vpwr_R_451 sky130_fd_sc_hd__decap_12
XDC_R_0_452 VGND VNB vpwr_R_452 vpwr_R_452 sky130_fd_sc_hd__decap_12
XDC_R_1_452 VGND VNB vpwr_R_452 vpwr_R_452 sky130_fd_sc_hd__decap_12
XDC_R_2_452 VGND VNB vpwr_R_452 vpwr_R_452 sky130_fd_sc_hd__decap_12
XDC_R_0_453 VGND VNB vpwr_R_453 vpwr_R_453 sky130_fd_sc_hd__decap_12
XDC_R_1_453 VGND VNB vpwr_R_453 vpwr_R_453 sky130_fd_sc_hd__decap_12
XDC_R_2_453 VGND VNB vpwr_R_453 vpwr_R_453 sky130_fd_sc_hd__decap_12
XDC_R_0_454 VGND VNB vpwr_R_454 vpwr_R_454 sky130_fd_sc_hd__decap_12
XDC_R_1_454 VGND VNB vpwr_R_454 vpwr_R_454 sky130_fd_sc_hd__decap_12
XDC_R_2_454 VGND VNB vpwr_R_454 vpwr_R_454 sky130_fd_sc_hd__decap_12
XDC_R_0_455 VGND VNB vpwr_R_455 vpwr_R_455 sky130_fd_sc_hd__decap_12
XDC_R_1_455 VGND VNB vpwr_R_455 vpwr_R_455 sky130_fd_sc_hd__decap_12
XDC_R_2_455 VGND VNB vpwr_R_455 vpwr_R_455 sky130_fd_sc_hd__decap_12
XDC_R_0_456 VGND VNB vpwr_R_456 vpwr_R_456 sky130_fd_sc_hd__decap_12
XDC_R_1_456 VGND VNB vpwr_R_456 vpwr_R_456 sky130_fd_sc_hd__decap_12
XDC_R_2_456 VGND VNB vpwr_R_456 vpwr_R_456 sky130_fd_sc_hd__decap_12
XDC_R_0_457 VGND VNB vpwr_R_457 vpwr_R_457 sky130_fd_sc_hd__decap_12
XDC_R_1_457 VGND VNB vpwr_R_457 vpwr_R_457 sky130_fd_sc_hd__decap_12
XDC_R_2_457 VGND VNB vpwr_R_457 vpwr_R_457 sky130_fd_sc_hd__decap_12
XDC_R_0_458 VGND VNB vpwr_R_458 vpwr_R_458 sky130_fd_sc_hd__decap_12
XDC_R_1_458 VGND VNB vpwr_R_458 vpwr_R_458 sky130_fd_sc_hd__decap_12
XDC_R_2_458 VGND VNB vpwr_R_458 vpwr_R_458 sky130_fd_sc_hd__decap_12
XDC_R_0_459 VGND VNB vpwr_R_459 vpwr_R_459 sky130_fd_sc_hd__decap_12
XDC_R_1_459 VGND VNB vpwr_R_459 vpwr_R_459 sky130_fd_sc_hd__decap_12
XDC_R_2_459 VGND VNB vpwr_R_459 vpwr_R_459 sky130_fd_sc_hd__decap_12
XDC_R_0_460 VGND VNB vpwr_R_460 vpwr_R_460 sky130_fd_sc_hd__decap_12
XDC_R_1_460 VGND VNB vpwr_R_460 vpwr_R_460 sky130_fd_sc_hd__decap_12
XDC_R_2_460 VGND VNB vpwr_R_460 vpwr_R_460 sky130_fd_sc_hd__decap_12
XDC_R_0_461 VGND VNB vpwr_R_461 vpwr_R_461 sky130_fd_sc_hd__decap_12
XDC_R_1_461 VGND VNB vpwr_R_461 vpwr_R_461 sky130_fd_sc_hd__decap_12
XDC_R_2_461 VGND VNB vpwr_R_461 vpwr_R_461 sky130_fd_sc_hd__decap_12
XDC_R_0_462 VGND VNB vpwr_R_462 vpwr_R_462 sky130_fd_sc_hd__decap_12
XDC_R_1_462 VGND VNB vpwr_R_462 vpwr_R_462 sky130_fd_sc_hd__decap_12
XDC_R_2_462 VGND VNB vpwr_R_462 vpwr_R_462 sky130_fd_sc_hd__decap_12
XDC_R_0_463 VGND VNB vpwr_R_463 vpwr_R_463 sky130_fd_sc_hd__decap_12
XDC_R_1_463 VGND VNB vpwr_R_463 vpwr_R_463 sky130_fd_sc_hd__decap_12
XDC_R_2_463 VGND VNB vpwr_R_463 vpwr_R_463 sky130_fd_sc_hd__decap_12
XDC_R_0_464 VGND VNB vpwr_R_464 vpwr_R_464 sky130_fd_sc_hd__decap_12
XDC_R_1_464 VGND VNB vpwr_R_464 vpwr_R_464 sky130_fd_sc_hd__decap_12
XDC_R_2_464 VGND VNB vpwr_R_464 vpwr_R_464 sky130_fd_sc_hd__decap_12
XDC_R_0_465 VGND VNB vpwr_R_465 vpwr_R_465 sky130_fd_sc_hd__decap_12
XDC_R_1_465 VGND VNB vpwr_R_465 vpwr_R_465 sky130_fd_sc_hd__decap_12
XDC_R_2_465 VGND VNB vpwr_R_465 vpwr_R_465 sky130_fd_sc_hd__decap_12
XDC_R_0_466 VGND VNB vpwr_R_466 vpwr_R_466 sky130_fd_sc_hd__decap_12
XDC_R_1_466 VGND VNB vpwr_R_466 vpwr_R_466 sky130_fd_sc_hd__decap_12
XDC_R_2_466 VGND VNB vpwr_R_466 vpwr_R_466 sky130_fd_sc_hd__decap_12
XDC_R_0_467 VGND VNB vpwr_R_467 vpwr_R_467 sky130_fd_sc_hd__decap_12
XDC_R_1_467 VGND VNB vpwr_R_467 vpwr_R_467 sky130_fd_sc_hd__decap_12
XDC_R_2_467 VGND VNB vpwr_R_467 vpwr_R_467 sky130_fd_sc_hd__decap_12
XDC_R_0_468 VGND VNB vpwr_R_468 vpwr_R_468 sky130_fd_sc_hd__decap_12
XDC_R_1_468 VGND VNB vpwr_R_468 vpwr_R_468 sky130_fd_sc_hd__decap_12
XDC_R_2_468 VGND VNB vpwr_R_468 vpwr_R_468 sky130_fd_sc_hd__decap_12
XDC_R_0_469 VGND VNB vpwr_R_469 vpwr_R_469 sky130_fd_sc_hd__decap_12
XDC_R_1_469 VGND VNB vpwr_R_469 vpwr_R_469 sky130_fd_sc_hd__decap_12
XDC_R_2_469 VGND VNB vpwr_R_469 vpwr_R_469 sky130_fd_sc_hd__decap_12
XDC_R_0_470 VGND VNB vpwr_R_470 vpwr_R_470 sky130_fd_sc_hd__decap_12
XDC_R_1_470 VGND VNB vpwr_R_470 vpwr_R_470 sky130_fd_sc_hd__decap_12
XDC_R_2_470 VGND VNB vpwr_R_470 vpwr_R_470 sky130_fd_sc_hd__decap_12
XDC_R_0_471 VGND VNB vpwr_R_471 vpwr_R_471 sky130_fd_sc_hd__decap_12
XDC_R_1_471 VGND VNB vpwr_R_471 vpwr_R_471 sky130_fd_sc_hd__decap_12
XDC_R_2_471 VGND VNB vpwr_R_471 vpwr_R_471 sky130_fd_sc_hd__decap_12
XDC_R_0_472 VGND VNB vpwr_R_472 vpwr_R_472 sky130_fd_sc_hd__decap_12
XDC_R_1_472 VGND VNB vpwr_R_472 vpwr_R_472 sky130_fd_sc_hd__decap_12
XDC_R_2_472 VGND VNB vpwr_R_472 vpwr_R_472 sky130_fd_sc_hd__decap_12
XDC_R_0_473 VGND VNB vpwr_R_473 vpwr_R_473 sky130_fd_sc_hd__decap_12
XDC_R_1_473 VGND VNB vpwr_R_473 vpwr_R_473 sky130_fd_sc_hd__decap_12
XDC_R_2_473 VGND VNB vpwr_R_473 vpwr_R_473 sky130_fd_sc_hd__decap_12
XDC_R_0_474 VGND VNB vpwr_R_474 vpwr_R_474 sky130_fd_sc_hd__decap_12
XDC_R_1_474 VGND VNB vpwr_R_474 vpwr_R_474 sky130_fd_sc_hd__decap_12
XDC_R_2_474 VGND VNB vpwr_R_474 vpwr_R_474 sky130_fd_sc_hd__decap_12
XDC_R_0_475 VGND VNB vpwr_R_475 vpwr_R_475 sky130_fd_sc_hd__decap_12
XDC_R_1_475 VGND VNB vpwr_R_475 vpwr_R_475 sky130_fd_sc_hd__decap_12
XDC_R_2_475 VGND VNB vpwr_R_475 vpwr_R_475 sky130_fd_sc_hd__decap_12
XDC_R_0_476 VGND VNB vpwr_R_476 vpwr_R_476 sky130_fd_sc_hd__decap_12
XDC_R_1_476 VGND VNB vpwr_R_476 vpwr_R_476 sky130_fd_sc_hd__decap_12
XDC_R_2_476 VGND VNB vpwr_R_476 vpwr_R_476 sky130_fd_sc_hd__decap_12
XDC_R_0_477 VGND VNB vpwr_R_477 vpwr_R_477 sky130_fd_sc_hd__decap_12
XDC_R_1_477 VGND VNB vpwr_R_477 vpwr_R_477 sky130_fd_sc_hd__decap_12
XDC_R_2_477 VGND VNB vpwr_R_477 vpwr_R_477 sky130_fd_sc_hd__decap_12
XDC_R_0_478 VGND VNB vpwr_R_478 vpwr_R_478 sky130_fd_sc_hd__decap_12
XDC_R_1_478 VGND VNB vpwr_R_478 vpwr_R_478 sky130_fd_sc_hd__decap_12
XDC_R_2_478 VGND VNB vpwr_R_478 vpwr_R_478 sky130_fd_sc_hd__decap_12
XDC_R_0_479 VGND VNB vpwr_R_479 vpwr_R_479 sky130_fd_sc_hd__decap_12
XDC_R_1_479 VGND VNB vpwr_R_479 vpwr_R_479 sky130_fd_sc_hd__decap_12
XDC_R_2_479 VGND VNB vpwr_R_479 vpwr_R_479 sky130_fd_sc_hd__decap_12
XDC_R_0_480 VGND VNB vpwr_R_480 vpwr_R_480 sky130_fd_sc_hd__decap_12
XDC_R_1_480 VGND VNB vpwr_R_480 vpwr_R_480 sky130_fd_sc_hd__decap_12
XDC_R_2_480 VGND VNB vpwr_R_480 vpwr_R_480 sky130_fd_sc_hd__decap_12
XDC_R_0_481 VGND VNB vpwr_R_481 vpwr_R_481 sky130_fd_sc_hd__decap_12
XDC_R_1_481 VGND VNB vpwr_R_481 vpwr_R_481 sky130_fd_sc_hd__decap_12
XDC_R_2_481 VGND VNB vpwr_R_481 vpwr_R_481 sky130_fd_sc_hd__decap_12
XDC_R_0_482 VGND VNB vpwr_R_482 vpwr_R_482 sky130_fd_sc_hd__decap_12
XDC_R_1_482 VGND VNB vpwr_R_482 vpwr_R_482 sky130_fd_sc_hd__decap_12
XDC_R_2_482 VGND VNB vpwr_R_482 vpwr_R_482 sky130_fd_sc_hd__decap_12
XDC_R_0_483 VGND VNB vpwr_R_483 vpwr_R_483 sky130_fd_sc_hd__decap_12
XDC_R_1_483 VGND VNB vpwr_R_483 vpwr_R_483 sky130_fd_sc_hd__decap_12
XDC_R_2_483 VGND VNB vpwr_R_483 vpwr_R_483 sky130_fd_sc_hd__decap_12
XDC_R_0_484 VGND VNB vpwr_R_484 vpwr_R_484 sky130_fd_sc_hd__decap_12
XDC_R_1_484 VGND VNB vpwr_R_484 vpwr_R_484 sky130_fd_sc_hd__decap_12
XDC_R_2_484 VGND VNB vpwr_R_484 vpwr_R_484 sky130_fd_sc_hd__decap_12
XDC_R_0_485 VGND VNB vpwr_R_485 vpwr_R_485 sky130_fd_sc_hd__decap_12
XDC_R_1_485 VGND VNB vpwr_R_485 vpwr_R_485 sky130_fd_sc_hd__decap_12
XDC_R_2_485 VGND VNB vpwr_R_485 vpwr_R_485 sky130_fd_sc_hd__decap_12
XDC_R_0_486 VGND VNB vpwr_R_486 vpwr_R_486 sky130_fd_sc_hd__decap_12
XDC_R_1_486 VGND VNB vpwr_R_486 vpwr_R_486 sky130_fd_sc_hd__decap_12
XDC_R_2_486 VGND VNB vpwr_R_486 vpwr_R_486 sky130_fd_sc_hd__decap_12
XDC_R_0_487 VGND VNB vpwr_R_487 vpwr_R_487 sky130_fd_sc_hd__decap_12
XDC_R_1_487 VGND VNB vpwr_R_487 vpwr_R_487 sky130_fd_sc_hd__decap_12
XDC_R_2_487 VGND VNB vpwr_R_487 vpwr_R_487 sky130_fd_sc_hd__decap_12
XDC_R_0_488 VGND VNB vpwr_R_488 vpwr_R_488 sky130_fd_sc_hd__decap_12
XDC_R_1_488 VGND VNB vpwr_R_488 vpwr_R_488 sky130_fd_sc_hd__decap_12
XDC_R_2_488 VGND VNB vpwr_R_488 vpwr_R_488 sky130_fd_sc_hd__decap_12
XDC_R_0_489 VGND VNB vpwr_R_489 vpwr_R_489 sky130_fd_sc_hd__decap_12
XDC_R_1_489 VGND VNB vpwr_R_489 vpwr_R_489 sky130_fd_sc_hd__decap_12
XDC_R_2_489 VGND VNB vpwr_R_489 vpwr_R_489 sky130_fd_sc_hd__decap_12
XDC_R_0_490 VGND VNB vpwr_R_490 vpwr_R_490 sky130_fd_sc_hd__decap_12
XDC_R_1_490 VGND VNB vpwr_R_490 vpwr_R_490 sky130_fd_sc_hd__decap_12
XDC_R_2_490 VGND VNB vpwr_R_490 vpwr_R_490 sky130_fd_sc_hd__decap_12
XDC_R_0_491 VGND VNB vpwr_R_491 vpwr_R_491 sky130_fd_sc_hd__decap_12
XDC_R_1_491 VGND VNB vpwr_R_491 vpwr_R_491 sky130_fd_sc_hd__decap_12
XDC_R_2_491 VGND VNB vpwr_R_491 vpwr_R_491 sky130_fd_sc_hd__decap_12
XDC_R_0_492 VGND VNB vpwr_R_492 vpwr_R_492 sky130_fd_sc_hd__decap_12
XDC_R_1_492 VGND VNB vpwr_R_492 vpwr_R_492 sky130_fd_sc_hd__decap_12
XDC_R_2_492 VGND VNB vpwr_R_492 vpwr_R_492 sky130_fd_sc_hd__decap_12
XDC_R_0_493 VGND VNB vpwr_R_493 vpwr_R_493 sky130_fd_sc_hd__decap_12
XDC_R_1_493 VGND VNB vpwr_R_493 vpwr_R_493 sky130_fd_sc_hd__decap_12
XDC_R_2_493 VGND VNB vpwr_R_493 vpwr_R_493 sky130_fd_sc_hd__decap_12
XDC_R_0_494 VGND VNB vpwr_R_494 vpwr_R_494 sky130_fd_sc_hd__decap_12
XDC_R_1_494 VGND VNB vpwr_R_494 vpwr_R_494 sky130_fd_sc_hd__decap_12
XDC_R_2_494 VGND VNB vpwr_R_494 vpwr_R_494 sky130_fd_sc_hd__decap_12
XDC_R_0_495 VGND VNB vpwr_R_495 vpwr_R_495 sky130_fd_sc_hd__decap_12
XDC_R_1_495 VGND VNB vpwr_R_495 vpwr_R_495 sky130_fd_sc_hd__decap_12
XDC_R_2_495 VGND VNB vpwr_R_495 vpwr_R_495 sky130_fd_sc_hd__decap_12
XDC_R_0_496 VGND VNB vpwr_R_496 vpwr_R_496 sky130_fd_sc_hd__decap_12
XDC_R_1_496 VGND VNB vpwr_R_496 vpwr_R_496 sky130_fd_sc_hd__decap_12
XDC_R_2_496 VGND VNB vpwr_R_496 vpwr_R_496 sky130_fd_sc_hd__decap_12
XDC_R_0_497 VGND VNB vpwr_R_497 vpwr_R_497 sky130_fd_sc_hd__decap_12
XDC_R_1_497 VGND VNB vpwr_R_497 vpwr_R_497 sky130_fd_sc_hd__decap_12
XDC_R_2_497 VGND VNB vpwr_R_497 vpwr_R_497 sky130_fd_sc_hd__decap_12
XDC_R_0_498 VGND VNB vpwr_R_498 vpwr_R_498 sky130_fd_sc_hd__decap_12
XDC_R_1_498 VGND VNB vpwr_R_498 vpwr_R_498 sky130_fd_sc_hd__decap_12
XDC_R_2_498 VGND VNB vpwr_R_498 vpwr_R_498 sky130_fd_sc_hd__decap_12
XDC_R_0_499 VGND VNB vpwr_R_499 vpwr_R_499 sky130_fd_sc_hd__decap_12
XDC_R_1_499 VGND VNB vpwr_R_499 vpwr_R_499 sky130_fd_sc_hd__decap_12
XDC_R_2_499 VGND VNB vpwr_R_499 vpwr_R_499 sky130_fd_sc_hd__decap_12
XDC_R_0_500 VGND VNB vpwr_R_500 vpwr_R_500 sky130_fd_sc_hd__decap_12
XDC_R_1_500 VGND VNB vpwr_R_500 vpwr_R_500 sky130_fd_sc_hd__decap_12
XDC_R_2_500 VGND VNB vpwr_R_500 vpwr_R_500 sky130_fd_sc_hd__decap_12
XDC_R_0_501 VGND VNB vpwr_R_501 vpwr_R_501 sky130_fd_sc_hd__decap_12
XDC_R_1_501 VGND VNB vpwr_R_501 vpwr_R_501 sky130_fd_sc_hd__decap_12
XDC_R_2_501 VGND VNB vpwr_R_501 vpwr_R_501 sky130_fd_sc_hd__decap_12
XDC_R_0_502 VGND VNB vpwr_R_502 vpwr_R_502 sky130_fd_sc_hd__decap_12
XDC_R_1_502 VGND VNB vpwr_R_502 vpwr_R_502 sky130_fd_sc_hd__decap_12
XDC_R_2_502 VGND VNB vpwr_R_502 vpwr_R_502 sky130_fd_sc_hd__decap_12
XDC_R_0_503 VGND VNB vpwr_R_503 vpwr_R_503 sky130_fd_sc_hd__decap_12
XDC_R_1_503 VGND VNB vpwr_R_503 vpwr_R_503 sky130_fd_sc_hd__decap_12
XDC_R_2_503 VGND VNB vpwr_R_503 vpwr_R_503 sky130_fd_sc_hd__decap_12
XDC_R_0_504 VGND VNB vpwr_R_504 vpwr_R_504 sky130_fd_sc_hd__decap_12
XDC_R_1_504 VGND VNB vpwr_R_504 vpwr_R_504 sky130_fd_sc_hd__decap_12
XDC_R_2_504 VGND VNB vpwr_R_504 vpwr_R_504 sky130_fd_sc_hd__decap_12
XDC_R_0_505 VGND VNB vpwr_R_505 vpwr_R_505 sky130_fd_sc_hd__decap_12
XDC_R_1_505 VGND VNB vpwr_R_505 vpwr_R_505 sky130_fd_sc_hd__decap_12
XDC_R_2_505 VGND VNB vpwr_R_505 vpwr_R_505 sky130_fd_sc_hd__decap_12
XDC_R_0_506 VGND VNB vpwr_R_506 vpwr_R_506 sky130_fd_sc_hd__decap_12
XDC_R_1_506 VGND VNB vpwr_R_506 vpwr_R_506 sky130_fd_sc_hd__decap_12
XDC_R_2_506 VGND VNB vpwr_R_506 vpwr_R_506 sky130_fd_sc_hd__decap_12
XDC_R_0_507 VGND VNB vpwr_R_507 vpwr_R_507 sky130_fd_sc_hd__decap_12
XDC_R_1_507 VGND VNB vpwr_R_507 vpwr_R_507 sky130_fd_sc_hd__decap_12
XDC_R_2_507 VGND VNB vpwr_R_507 vpwr_R_507 sky130_fd_sc_hd__decap_12
XDC_R_0_508 VGND VNB vpwr_R_508 vpwr_R_508 sky130_fd_sc_hd__decap_12
XDC_R_1_508 VGND VNB vpwr_R_508 vpwr_R_508 sky130_fd_sc_hd__decap_12
XDC_R_2_508 VGND VNB vpwr_R_508 vpwr_R_508 sky130_fd_sc_hd__decap_12
XDC_R_0_509 VGND VNB vpwr_R_509 vpwr_R_509 sky130_fd_sc_hd__decap_12
XDC_R_1_509 VGND VNB vpwr_R_509 vpwr_R_509 sky130_fd_sc_hd__decap_12
XDC_R_2_509 VGND VNB vpwr_R_509 vpwr_R_509 sky130_fd_sc_hd__decap_12
XDC_R_0_510 VGND VNB vpwr_R_510 vpwr_R_510 sky130_fd_sc_hd__decap_12
XDC_R_1_510 VGND VNB vpwr_R_510 vpwr_R_510 sky130_fd_sc_hd__decap_12
XDC_R_2_510 VGND VNB vpwr_R_510 vpwr_R_510 sky130_fd_sc_hd__decap_12
XDC_R_0_511 VGND VNB vpwr_R_511 vpwr_R_511 sky130_fd_sc_hd__decap_12
XDC_R_1_511 VGND VNB vpwr_R_511 vpwr_R_511 sky130_fd_sc_hd__decap_12
XDC_R_2_511 VGND VNB vpwr_R_511 vpwr_R_511 sky130_fd_sc_hd__decap_12
XDC_R_0_512 VGND VNB vpwr_R_512 vpwr_R_512 sky130_fd_sc_hd__decap_12
XDC_R_1_512 VGND VNB vpwr_R_512 vpwr_R_512 sky130_fd_sc_hd__decap_12
XDC_R_2_512 VGND VNB vpwr_R_512 vpwr_R_512 sky130_fd_sc_hd__decap_12
XDC_R_0_513 VGND VNB vpwr_R_513 vpwr_R_513 sky130_fd_sc_hd__decap_12
XDC_R_1_513 VGND VNB vpwr_R_513 vpwr_R_513 sky130_fd_sc_hd__decap_12
XDC_R_2_513 VGND VNB vpwr_R_513 vpwr_R_513 sky130_fd_sc_hd__decap_12
XDC_R_0_514 VGND VNB vpwr_R_514 vpwr_R_514 sky130_fd_sc_hd__decap_12
XDC_R_1_514 VGND VNB vpwr_R_514 vpwr_R_514 sky130_fd_sc_hd__decap_12
XDC_R_2_514 VGND VNB vpwr_R_514 vpwr_R_514 sky130_fd_sc_hd__decap_12
XDC_R_0_515 VGND VNB vpwr_R_515 vpwr_R_515 sky130_fd_sc_hd__decap_12
XDC_R_1_515 VGND VNB vpwr_R_515 vpwr_R_515 sky130_fd_sc_hd__decap_12
XDC_R_2_515 VGND VNB vpwr_R_515 vpwr_R_515 sky130_fd_sc_hd__decap_12
XDC_R_0_516 VGND VNB vpwr_R_516 vpwr_R_516 sky130_fd_sc_hd__decap_12
XDC_R_1_516 VGND VNB vpwr_R_516 vpwr_R_516 sky130_fd_sc_hd__decap_12
XDC_R_2_516 VGND VNB vpwr_R_516 vpwr_R_516 sky130_fd_sc_hd__decap_12
XDC_R_0_517 VGND VNB vpwr_R_517 vpwr_R_517 sky130_fd_sc_hd__decap_12
XDC_R_1_517 VGND VNB vpwr_R_517 vpwr_R_517 sky130_fd_sc_hd__decap_12
XDC_R_2_517 VGND VNB vpwr_R_517 vpwr_R_517 sky130_fd_sc_hd__decap_12
XDC_R_0_518 VGND VNB vpwr_R_518 vpwr_R_518 sky130_fd_sc_hd__decap_12
XDC_R_1_518 VGND VNB vpwr_R_518 vpwr_R_518 sky130_fd_sc_hd__decap_12
XDC_R_2_518 VGND VNB vpwr_R_518 vpwr_R_518 sky130_fd_sc_hd__decap_12
XDC_R_0_519 VGND VNB vpwr_R_519 vpwr_R_519 sky130_fd_sc_hd__decap_12
XDC_R_1_519 VGND VNB vpwr_R_519 vpwr_R_519 sky130_fd_sc_hd__decap_12
XDC_R_2_519 VGND VNB vpwr_R_519 vpwr_R_519 sky130_fd_sc_hd__decap_12
XDC_R_0_520 VGND VNB vpwr_R_520 vpwr_R_520 sky130_fd_sc_hd__decap_12
XDC_R_1_520 VGND VNB vpwr_R_520 vpwr_R_520 sky130_fd_sc_hd__decap_12
XDC_R_2_520 VGND VNB vpwr_R_520 vpwr_R_520 sky130_fd_sc_hd__decap_12
XDC_R_0_521 VGND VNB vpwr_R_521 vpwr_R_521 sky130_fd_sc_hd__decap_12
XDC_R_1_521 VGND VNB vpwr_R_521 vpwr_R_521 sky130_fd_sc_hd__decap_12
XDC_R_2_521 VGND VNB vpwr_R_521 vpwr_R_521 sky130_fd_sc_hd__decap_12
XDC_R_0_522 VGND VNB vpwr_R_522 vpwr_R_522 sky130_fd_sc_hd__decap_12
XDC_R_1_522 VGND VNB vpwr_R_522 vpwr_R_522 sky130_fd_sc_hd__decap_12
XDC_R_2_522 VGND VNB vpwr_R_522 vpwr_R_522 sky130_fd_sc_hd__decap_12
XDC_R_0_523 VGND VNB vpwr_R_523 vpwr_R_523 sky130_fd_sc_hd__decap_12
XDC_R_1_523 VGND VNB vpwr_R_523 vpwr_R_523 sky130_fd_sc_hd__decap_12
XDC_R_2_523 VGND VNB vpwr_R_523 vpwr_R_523 sky130_fd_sc_hd__decap_12
XDC_R_0_524 VGND VNB vpwr_R_524 vpwr_R_524 sky130_fd_sc_hd__decap_12
XDC_R_1_524 VGND VNB vpwr_R_524 vpwr_R_524 sky130_fd_sc_hd__decap_12
XDC_R_2_524 VGND VNB vpwr_R_524 vpwr_R_524 sky130_fd_sc_hd__decap_12
XDC_R_0_525 VGND VNB vpwr_R_525 vpwr_R_525 sky130_fd_sc_hd__decap_12
XDC_R_1_525 VGND VNB vpwr_R_525 vpwr_R_525 sky130_fd_sc_hd__decap_12
XDC_R_2_525 VGND VNB vpwr_R_525 vpwr_R_525 sky130_fd_sc_hd__decap_12
XDC_R_0_526 VGND VNB vpwr_R_526 vpwr_R_526 sky130_fd_sc_hd__decap_12
XDC_R_1_526 VGND VNB vpwr_R_526 vpwr_R_526 sky130_fd_sc_hd__decap_12
XDC_R_2_526 VGND VNB vpwr_R_526 vpwr_R_526 sky130_fd_sc_hd__decap_12
XDC_R_0_527 VGND VNB vpwr_R_527 vpwr_R_527 sky130_fd_sc_hd__decap_12
XDC_R_1_527 VGND VNB vpwr_R_527 vpwr_R_527 sky130_fd_sc_hd__decap_12
XDC_R_2_527 VGND VNB vpwr_R_527 vpwr_R_527 sky130_fd_sc_hd__decap_12
XDC_R_0_528 VGND VNB vpwr_R_528 vpwr_R_528 sky130_fd_sc_hd__decap_12
XDC_R_1_528 VGND VNB vpwr_R_528 vpwr_R_528 sky130_fd_sc_hd__decap_12
XDC_R_2_528 VGND VNB vpwr_R_528 vpwr_R_528 sky130_fd_sc_hd__decap_12
XDC_R_0_529 VGND VNB vpwr_R_529 vpwr_R_529 sky130_fd_sc_hd__decap_12
XDC_R_1_529 VGND VNB vpwr_R_529 vpwr_R_529 sky130_fd_sc_hd__decap_12
XDC_R_2_529 VGND VNB vpwr_R_529 vpwr_R_529 sky130_fd_sc_hd__decap_12
XDC_R_0_530 VGND VNB vpwr_R_530 vpwr_R_530 sky130_fd_sc_hd__decap_12
XDC_R_1_530 VGND VNB vpwr_R_530 vpwr_R_530 sky130_fd_sc_hd__decap_12
XDC_R_2_530 VGND VNB vpwr_R_530 vpwr_R_530 sky130_fd_sc_hd__decap_12
XDC_R_0_531 VGND VNB vpwr_R_531 vpwr_R_531 sky130_fd_sc_hd__decap_12
XDC_R_1_531 VGND VNB vpwr_R_531 vpwr_R_531 sky130_fd_sc_hd__decap_12
XDC_R_2_531 VGND VNB vpwr_R_531 vpwr_R_531 sky130_fd_sc_hd__decap_12
XDC_R_0_532 VGND VNB vpwr_R_532 vpwr_R_532 sky130_fd_sc_hd__decap_12
XDC_R_1_532 VGND VNB vpwr_R_532 vpwr_R_532 sky130_fd_sc_hd__decap_12
XDC_R_2_532 VGND VNB vpwr_R_532 vpwr_R_532 sky130_fd_sc_hd__decap_12
XDC_R_0_533 VGND VNB vpwr_R_533 vpwr_R_533 sky130_fd_sc_hd__decap_12
XDC_R_1_533 VGND VNB vpwr_R_533 vpwr_R_533 sky130_fd_sc_hd__decap_12
XDC_R_2_533 VGND VNB vpwr_R_533 vpwr_R_533 sky130_fd_sc_hd__decap_12
XDC_R_0_534 VGND VNB vpwr_R_534 vpwr_R_534 sky130_fd_sc_hd__decap_12
XDC_R_1_534 VGND VNB vpwr_R_534 vpwr_R_534 sky130_fd_sc_hd__decap_12
XDC_R_2_534 VGND VNB vpwr_R_534 vpwr_R_534 sky130_fd_sc_hd__decap_12
XDC_R_0_535 VGND VNB vpwr_R_535 vpwr_R_535 sky130_fd_sc_hd__decap_12
XDC_R_1_535 VGND VNB vpwr_R_535 vpwr_R_535 sky130_fd_sc_hd__decap_12
XDC_R_2_535 VGND VNB vpwr_R_535 vpwr_R_535 sky130_fd_sc_hd__decap_12
XDC_R_0_536 VGND VNB vpwr_R_536 vpwr_R_536 sky130_fd_sc_hd__decap_12
XDC_R_1_536 VGND VNB vpwr_R_536 vpwr_R_536 sky130_fd_sc_hd__decap_12
XDC_R_2_536 VGND VNB vpwr_R_536 vpwr_R_536 sky130_fd_sc_hd__decap_12
XDC_R_0_537 VGND VNB vpwr_R_537 vpwr_R_537 sky130_fd_sc_hd__decap_12
XDC_R_1_537 VGND VNB vpwr_R_537 vpwr_R_537 sky130_fd_sc_hd__decap_12
XDC_R_2_537 VGND VNB vpwr_R_537 vpwr_R_537 sky130_fd_sc_hd__decap_12
XDC_R_0_538 VGND VNB vpwr_R_538 vpwr_R_538 sky130_fd_sc_hd__decap_12
XDC_R_1_538 VGND VNB vpwr_R_538 vpwr_R_538 sky130_fd_sc_hd__decap_12
XDC_R_2_538 VGND VNB vpwr_R_538 vpwr_R_538 sky130_fd_sc_hd__decap_12
XDC_R_0_539 VGND VNB vpwr_R_539 vpwr_R_539 sky130_fd_sc_hd__decap_12
XDC_R_1_539 VGND VNB vpwr_R_539 vpwr_R_539 sky130_fd_sc_hd__decap_12
XDC_R_2_539 VGND VNB vpwr_R_539 vpwr_R_539 sky130_fd_sc_hd__decap_12
XDC_R_0_540 VGND VNB vpwr_R_540 vpwr_R_540 sky130_fd_sc_hd__decap_12
XDC_R_1_540 VGND VNB vpwr_R_540 vpwr_R_540 sky130_fd_sc_hd__decap_12
XDC_R_2_540 VGND VNB vpwr_R_540 vpwr_R_540 sky130_fd_sc_hd__decap_12
XDC_R_0_541 VGND VNB vpwr_R_541 vpwr_R_541 sky130_fd_sc_hd__decap_12
XDC_R_1_541 VGND VNB vpwr_R_541 vpwr_R_541 sky130_fd_sc_hd__decap_12
XDC_R_2_541 VGND VNB vpwr_R_541 vpwr_R_541 sky130_fd_sc_hd__decap_12
XDC_R_0_542 VGND VNB vpwr_R_542 vpwr_R_542 sky130_fd_sc_hd__decap_12
XDC_R_1_542 VGND VNB vpwr_R_542 vpwr_R_542 sky130_fd_sc_hd__decap_12
XDC_R_2_542 VGND VNB vpwr_R_542 vpwr_R_542 sky130_fd_sc_hd__decap_12
XDC_R_0_543 VGND VNB vpwr_R_543 vpwr_R_543 sky130_fd_sc_hd__decap_12
XDC_R_1_543 VGND VNB vpwr_R_543 vpwr_R_543 sky130_fd_sc_hd__decap_12
XDC_R_2_543 VGND VNB vpwr_R_543 vpwr_R_543 sky130_fd_sc_hd__decap_12

VC_0  clk_0  VGND pulse 0 1.8 1.34n 1n 1n 48n 100n
VC_1  clk_1  VGND pulse 0 1.8 0.99n 1n 1n 48n 100n
VC_2  clk_2  VGND pulse 0 1.8 1.21n 1n 1n 48n 100n
VC_3  clk_3  VGND pulse 0 1.8  0.4n 1n 1n 48n 100n
VC_4  clk_4  VGND pulse 0 1.8 0.01n 1n 1n 48n 100n
VC_5  clk_5  VGND pulse 0 1.8 0.82n 1n 1n 48n 100n
VC_6  clk_6  VGND pulse 0 1.8 0.31n 1n 1n 48n 100n
VC_7  clk_7  VGND pulse 0 1.8 1.06n 1n 1n 48n 100n
VC_8  clk_8  VGND pulse 0 1.8 1.27n 1n 1n 48n 100n
VC_9  clk_9  VGND pulse 0 1.8 0.18n 1n 1n 48n 100n
VC_10 clk_10 VGND pulse 0 1.8 0.39n 1n 1n 48n 100n
VC_11 clk_11 VGND pulse 0 1.8 1.19n 1n 1n 48n 100n
VC_12 clk_12 VGND pulse 0 1.8  1.3n 1n 1n 48n 100n
VC_13 clk_13 VGND pulse 0 1.8 0.07n 1n 1n 48n 100n
VC_14 clk_14 VGND pulse 0 1.8 1.24n 1n 1n 48n 100n
VC_15 clk_15 VGND pulse 0 1.8 1.14n 1n 1n 48n 100n
VC_16 clk_16 VGND pulse 0 1.8 1.18n 1n 1n 48n 100n
VC_17 clk_17 VGND pulse 0 1.8 1.29n 1n 1n 48n 100n
VC_18 clk_18 VGND pulse 0 1.8 0.71n 1n 1n 48n 100n
VC_19 clk_19 VGND pulse 0 1.8 0.82n 1n 1n 48n 100n
VC_20 clk_20 VGND pulse 0 1.8  1.4n 1n 1n 48n 100n
VC_21 clk_21 VGND pulse 0 1.8 1.07n 1n 1n 48n 100n
VC_22 clk_22 VGND pulse 0 1.8 1.17n 1n 1n 48n 100n
VC_23 clk_23 VGND pulse 0 1.8 0.36n 1n 1n 48n 100n
VC_24 clk_24 VGND pulse 0 1.8 0.21n 1n 1n 48n 100n
VC_25 clk_25 VGND pulse 0 1.8 0.87n 1n 1n 48n 100n
VC_26 clk_26 VGND pulse 0 1.8 0.78n 1n 1n 48n 100n
VC_27 clk_27 VGND pulse 0 1.8  1.1n 1n 1n 48n 100n
VC_28 clk_28 VGND pulse 0 1.8 0.37n 1n 1n 48n 100n
VC_29 clk_29 VGND pulse 0 1.8 1.16n 1n 1n 48n 100n
VC_30 clk_30 VGND pulse 0 1.8 1.35n 1n 1n 48n 100n
VC_31 clk_31 VGND pulse 0 1.8 0.43n 1n 1n 48n 100n

x1_0  clk_0  VGND VNB vpwr_R_0  vpwr_R_0  co_0  sky130_fd_sc_hd__clkbuf_1
x1_1  clk_1  VGND VNB vpwr_R_10 vpwr_R_10 co_1  sky130_fd_sc_hd__clkbuf_1
x1_2  clk_2  VGND VNB vpwr_R_22 vpwr_R_22 co_2  sky130_fd_sc_hd__clkbuf_1
x1_3  clk_3  VGND VNB vpwr_R_31 vpwr_R_31 co_3  sky130_fd_sc_hd__clkbuf_1
x1_4  clk_4  VGND VNB vpwr_R_40 vpwr_R_40 co_4  sky130_fd_sc_hd__clkbuf_1
x1_5  clk_5  VGND VNB vpwr_R_49 vpwr_R_49 co_5  sky130_fd_sc_hd__clkbuf_1
x1_6  clk_6  VGND VNB vpwr_R_62 vpwr_R_62 co_6  sky130_fd_sc_hd__clkbuf_1
x1_7  clk_7  VGND VNB vpwr_R_73 vpwr_R_73 co_7  sky130_fd_sc_hd__clkbuf_1
x1_8  clk_8  VGND VNB vpwr_R_89 vpwr_R_89 co_8  sky130_fd_sc_hd__clkbuf_1
x1_9  clk_9  VGND VNB vpwr_R_94 vpwr_R_94 co_9  sky130_fd_sc_hd__clkbuf_1
x1_10 clk_10 VGND VNB vpwr_R_100 vpwr_R_100 co_10 sky130_fd_sc_hd__clkbuf_1
x1_11 clk_11 VGND VNB vpwr_R_108 vpwr_R_108 co_11 sky130_fd_sc_hd__clkbuf_1
x1_12 clk_12 VGND VNB vpwr_R_117 vpwr_R_117 co_12 sky130_fd_sc_hd__clkbuf_1
x1_13 clk_13 VGND VNB vpwr_R_123 vpwr_R_123 co_13 sky130_fd_sc_hd__clkbuf_1
x1_14 clk_14 VGND VNB vpwr_R_131 vpwr_R_131 co_14 sky130_fd_sc_hd__clkbuf_1
x1_15 clk_15 VGND VNB vpwr_R_137 vpwr_R_137 co_15 sky130_fd_sc_hd__clkbuf_1
x1_16 clk_16 VGND VNB vpwr_R_145 vpwr_R_145 co_16 sky130_fd_sc_hd__clkbuf_1
x1_17 clk_17 VGND VNB vpwr_R_157 vpwr_R_157 co_17 sky130_fd_sc_hd__clkbuf_1
x1_18 clk_18 VGND VNB vpwr_R_172 vpwr_R_172 co_18 sky130_fd_sc_hd__clkbuf_1
x1_19 clk_19 VGND VNB vpwr_R_186 vpwr_R_186 co_19 sky130_fd_sc_hd__clkbuf_1
x1_20 clk_20 VGND VNB vpwr_R_195 vpwr_R_195 co_20 sky130_fd_sc_hd__clkbuf_1
x1_21 clk_21 VGND VNB vpwr_R_211 vpwr_R_211 co_21 sky130_fd_sc_hd__clkbuf_1
x1_22 clk_22 VGND VNB vpwr_R_225 vpwr_R_225 co_22 sky130_fd_sc_hd__clkbuf_1
x1_23 clk_23 VGND VNB vpwr_R_236 vpwr_R_236 co_23 sky130_fd_sc_hd__clkbuf_1
x1_24 clk_24 VGND VNB vpwr_R_253 vpwr_R_253 co_24 sky130_fd_sc_hd__clkbuf_1
x1_25 clk_25 VGND VNB vpwr_R_265 vpwr_R_265 co_25 sky130_fd_sc_hd__clkbuf_1
x1_26 clk_26 VGND VNB vpwr_R_278 vpwr_R_278 co_26 sky130_fd_sc_hd__clkbuf_1
x1_27 clk_27 VGND VNB vpwr_R_289 vpwr_R_289 co_27 sky130_fd_sc_hd__clkbuf_1
x1_28 clk_28 VGND VNB vpwr_R_299 vpwr_R_299 co_28 sky130_fd_sc_hd__clkbuf_1
x1_29 clk_29 VGND VNB vpwr_R_313 vpwr_R_313 co_29 sky130_fd_sc_hd__clkbuf_1
x1_30 clk_30 VGND VNB vpwr_R_327 vpwr_R_327 co_30 sky130_fd_sc_hd__clkbuf_1
x1_31 clk_31 VGND VNB vpwr_R_336 vpwr_R_336 co_31 sky130_fd_sc_hd__clkbuf_1

R_0  co_0  co_1  ${R_LOAD}
R_1  co_1  co_2  ${R_LOAD}
R_2  co_2  co_3  ${R_LOAD}
R_3  co_3  co_4  ${R_LOAD}
R_4  co_4  co_5  ${R_LOAD}
R_5  co_5  co_6  ${R_LOAD}
R_6  co_6  co_7  ${R_LOAD}
R_7  co_7  co_8  ${R_LOAD}
R_8  co_8  co_9  ${R_LOAD}
R_9  co_9  co_10 ${R_LOAD}
R_10 co_10 co_11 ${R_LOAD}
R_11 co_11 co_12 ${R_LOAD}
R_12 co_12 co_13 ${R_LOAD}
R_13 co_13 co_14 ${R_LOAD}
R_14 co_14 co_15 ${R_LOAD}
R_15 co_15 co_16 ${R_LOAD}
R_16 co_16 co_17 ${R_LOAD}
R_17 co_17 co_18 ${R_LOAD}
R_18 co_18 co_19 ${R_LOAD}
R_19 co_19 co_20 ${R_LOAD}
R_20 co_20 co_21 ${R_LOAD}
R_21 co_21 co_22 ${R_LOAD}
R_22 co_22 co_23 ${R_LOAD}
R_23 co_23 co_24 ${R_LOAD}
R_24 co_24 co_25 ${R_LOAD}
R_25 co_25 co_26 ${R_LOAD}
R_26 co_26 co_27 ${R_LOAD}
R_27 co_27 co_28 ${R_LOAD}
R_28 co_28 co_29 ${R_LOAD}
R_29 co_29 co_30 ${R_LOAD}
R_30 co_30 co_31 ${R_LOAD}
R_31 co_31 co_32 ${R_LOAD}

x_buf1_buf16_intcon_0_0  co_0 co_i_0_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_0_1  co_0 co_i_0_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_0_2  co_0 co_i_0_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_0_3  co_0 co_i_0_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_0_4  co_0 co_i_0_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_0_5  co_0 co_i_0_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_0_6  co_0 co_i_0_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_0_7  co_0 co_i_0_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_0_8  co_0 co_i_0_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_0  co_1 co_i_1_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_1  co_1 co_i_1_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_2  co_1 co_i_1_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_3  co_1 co_i_1_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_4  co_1 co_i_1_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_5  co_1 co_i_1_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_6  co_1 co_i_1_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_7  co_1 co_i_1_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_8  co_1 co_i_1_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_9  co_1 co_i_1_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_1_10 co_1 co_i_1_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_2_0  co_2 co_i_2_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_2_1  co_2 co_i_2_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_2_2  co_2 co_i_2_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_2_3  co_2 co_i_2_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_2_4  co_2 co_i_2_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_2_5  co_2 co_i_2_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_2_6  co_2 co_i_2_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_2_7  co_2 co_i_2_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_3_0  co_3 co_i_3_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_3_1  co_3 co_i_3_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_3_2  co_3 co_i_3_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_3_3  co_3 co_i_3_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_3_4  co_3 co_i_3_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_3_5  co_3 co_i_3_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_3_6  co_3 co_i_3_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_3_7  co_3 co_i_3_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_4_0  co_4 co_i_4_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_4_1  co_4 co_i_4_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_4_2  co_4 co_i_4_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_4_3  co_4 co_i_4_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_4_4  co_4 co_i_4_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_4_5  co_4 co_i_4_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_4_6  co_4 co_i_4_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_4_7  co_4 co_i_4_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_0  co_5 co_i_5_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_1  co_5 co_i_5_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_2  co_5 co_i_5_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_3  co_5 co_i_5_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_4  co_5 co_i_5_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_5  co_5 co_i_5_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_6  co_5 co_i_5_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_7  co_5 co_i_5_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_8  co_5 co_i_5_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_9  co_5 co_i_5_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_10 co_5 co_i_5_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_5_11 co_5 co_i_5_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_0  co_6 co_i_6_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_1  co_6 co_i_6_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_2  co_6 co_i_6_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_3  co_6 co_i_6_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_4  co_6 co_i_6_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_5  co_6 co_i_6_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_6  co_6 co_i_6_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_7  co_6 co_i_6_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_8  co_6 co_i_6_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_6_9  co_6 co_i_6_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_0  co_7 co_i_7_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_1  co_7 co_i_7_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_2  co_7 co_i_7_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_3  co_7 co_i_7_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_4  co_7 co_i_7_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_5  co_7 co_i_7_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_6  co_7 co_i_7_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_7  co_7 co_i_7_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_8  co_7 co_i_7_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_9  co_7 co_i_7_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_10 co_7 co_i_7_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_11 co_7 co_i_7_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_12 co_7 co_i_7_12 VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_13 co_7 co_i_7_13 VGND int_con C=8F R=120
x_buf1_buf16_intcon_7_14 co_7 co_i_7_14 VGND int_con C=8F R=120
x_buf1_buf16_intcon_8_0  co_8 co_i_8_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_8_1  co_8 co_i_8_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_8_2  co_8 co_i_8_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_8_3  co_8 co_i_8_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_9_0  co_9 co_i_9_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_9_1  co_9 co_i_9_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_9_2  co_9 co_i_9_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_9_3  co_9 co_i_9_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_9_4  co_9 co_i_9_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_10_0  co_10 co_i_10_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_10_1  co_10 co_i_10_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_10_2  co_10 co_i_10_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_10_3  co_10 co_i_10_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_10_4  co_10 co_i_10_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_10_5  co_10 co_i_10_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_10_6  co_10 co_i_10_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_11_0  co_11 co_i_11_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_11_1  co_11 co_i_11_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_11_2  co_11 co_i_11_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_11_3  co_11 co_i_11_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_11_4  co_11 co_i_11_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_11_5  co_11 co_i_11_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_11_6  co_11 co_i_11_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_11_7  co_11 co_i_11_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_12_0  co_12 co_i_12_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_12_1  co_12 co_i_12_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_12_2  co_12 co_i_12_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_12_3  co_12 co_i_12_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_12_4  co_12 co_i_12_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_13_0  co_13 co_i_13_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_13_1  co_13 co_i_13_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_13_2  co_13 co_i_13_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_13_3  co_13 co_i_13_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_13_4  co_13 co_i_13_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_13_5  co_13 co_i_13_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_13_6  co_13 co_i_13_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_14_0  co_14 co_i_14_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_14_1  co_14 co_i_14_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_14_2  co_14 co_i_14_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_14_3  co_14 co_i_14_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_14_4  co_14 co_i_14_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_15_0  co_15 co_i_15_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_15_1  co_15 co_i_15_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_15_2  co_15 co_i_15_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_15_3  co_15 co_i_15_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_15_4  co_15 co_i_15_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_15_5  co_15 co_i_15_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_15_6  co_15 co_i_15_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_0  co_16 co_i_16_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_1  co_16 co_i_16_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_2  co_16 co_i_16_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_3  co_16 co_i_16_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_4  co_16 co_i_16_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_5  co_16 co_i_16_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_6  co_16 co_i_16_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_7  co_16 co_i_16_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_8  co_16 co_i_16_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_9  co_16 co_i_16_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_16_10 co_16 co_i_16_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_0  co_17 co_i_17_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_1  co_17 co_i_17_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_2  co_17 co_i_17_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_3  co_17 co_i_17_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_4  co_17 co_i_17_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_5  co_17 co_i_17_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_6  co_17 co_i_17_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_7  co_17 co_i_17_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_8  co_17 co_i_17_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_9  co_17 co_i_17_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_10 co_17 co_i_17_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_11 co_17 co_i_17_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_12 co_17 co_i_17_12 VGND int_con C=8F R=120
x_buf1_buf16_intcon_17_13 co_17 co_i_17_13 VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_0  co_18 co_i_18_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_1  co_18 co_i_18_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_2  co_18 co_i_18_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_3  co_18 co_i_18_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_4  co_18 co_i_18_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_5  co_18 co_i_18_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_6  co_18 co_i_18_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_7  co_18 co_i_18_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_8  co_18 co_i_18_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_9  co_18 co_i_18_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_10 co_18 co_i_18_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_11 co_18 co_i_18_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_18_12 co_18 co_i_18_12 VGND int_con C=8F R=120
x_buf1_buf16_intcon_19_0  co_19 co_i_19_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_19_1  co_19 co_i_19_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_19_2  co_19 co_i_19_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_19_3  co_19 co_i_19_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_19_4  co_19 co_i_19_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_19_5  co_19 co_i_19_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_19_6  co_19 co_i_19_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_19_7  co_19 co_i_19_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_0  co_20 co_i_20_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_1  co_20 co_i_20_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_2  co_20 co_i_20_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_3  co_20 co_i_20_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_4  co_20 co_i_20_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_5  co_20 co_i_20_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_6  co_20 co_i_20_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_7  co_20 co_i_20_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_8  co_20 co_i_20_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_9  co_20 co_i_20_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_10 co_20 co_i_20_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_11 co_20 co_i_20_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_12 co_20 co_i_20_12 VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_13 co_20 co_i_20_13 VGND int_con C=8F R=120
x_buf1_buf16_intcon_20_14 co_20 co_i_20_14 VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_0  co_21 co_i_21_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_1  co_21 co_i_21_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_2  co_21 co_i_21_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_3  co_21 co_i_21_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_4  co_21 co_i_21_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_5  co_21 co_i_21_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_6  co_21 co_i_21_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_7  co_21 co_i_21_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_8  co_21 co_i_21_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_9  co_21 co_i_21_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_10 co_21 co_i_21_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_11 co_21 co_i_21_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_21_12 co_21 co_i_21_12 VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_0  co_22 co_i_22_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_1  co_22 co_i_22_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_2  co_22 co_i_22_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_3  co_22 co_i_22_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_4  co_22 co_i_22_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_5  co_22 co_i_22_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_6  co_22 co_i_22_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_7  co_22 co_i_22_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_8  co_22 co_i_22_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_22_9  co_22 co_i_22_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_0  co_23 co_i_23_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_1  co_23 co_i_23_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_2  co_23 co_i_23_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_3  co_23 co_i_23_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_4  co_23 co_i_23_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_5  co_23 co_i_23_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_6  co_23 co_i_23_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_7  co_23 co_i_23_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_8  co_23 co_i_23_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_9  co_23 co_i_23_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_10 co_23 co_i_23_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_11 co_23 co_i_23_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_12 co_23 co_i_23_12 VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_13 co_23 co_i_23_13 VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_14 co_23 co_i_23_14 VGND int_con C=8F R=120
x_buf1_buf16_intcon_23_15 co_23 co_i_23_15 VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_0  co_24 co_i_24_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_1  co_24 co_i_24_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_2  co_24 co_i_24_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_3  co_24 co_i_24_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_4  co_24 co_i_24_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_5  co_24 co_i_24_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_6  co_24 co_i_24_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_7  co_24 co_i_24_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_8  co_24 co_i_24_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_9  co_24 co_i_24_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_24_10 co_24 co_i_24_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_0  co_25 co_i_25_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_1  co_25 co_i_25_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_2  co_25 co_i_25_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_3  co_25 co_i_25_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_4  co_25 co_i_25_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_5  co_25 co_i_25_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_6  co_25 co_i_25_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_7  co_25 co_i_25_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_8  co_25 co_i_25_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_9  co_25 co_i_25_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_10 co_25 co_i_25_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_25_11 co_25 co_i_25_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_0  co_26 co_i_26_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_1  co_26 co_i_26_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_2  co_26 co_i_26_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_3  co_26 co_i_26_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_4  co_26 co_i_26_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_5  co_26 co_i_26_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_6  co_26 co_i_26_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_7  co_26 co_i_26_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_8  co_26 co_i_26_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_26_9  co_26 co_i_26_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_0  co_27 co_i_27_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_1  co_27 co_i_27_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_2  co_27 co_i_27_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_3  co_27 co_i_27_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_4  co_27 co_i_27_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_5  co_27 co_i_27_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_6  co_27 co_i_27_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_7  co_27 co_i_27_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_27_8  co_27 co_i_27_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_0  co_28 co_i_28_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_1  co_28 co_i_28_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_2  co_28 co_i_28_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_3  co_28 co_i_28_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_4  co_28 co_i_28_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_5  co_28 co_i_28_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_6  co_28 co_i_28_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_7  co_28 co_i_28_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_8  co_28 co_i_28_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_9  co_28 co_i_28_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_10 co_28 co_i_28_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_11 co_28 co_i_28_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_28_12 co_28 co_i_28_12 VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_0  co_29 co_i_29_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_1  co_29 co_i_29_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_2  co_29 co_i_29_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_3  co_29 co_i_29_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_4  co_29 co_i_29_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_5  co_29 co_i_29_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_6  co_29 co_i_29_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_7  co_29 co_i_29_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_8  co_29 co_i_29_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_9  co_29 co_i_29_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_10 co_29 co_i_29_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_11 co_29 co_i_29_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_29_12 co_29 co_i_29_12 VGND int_con C=8F R=120
x_buf1_buf16_intcon_30_0  co_30 co_i_30_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_30_1  co_30 co_i_30_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_30_2  co_30 co_i_30_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_30_3  co_30 co_i_30_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_30_4  co_30 co_i_30_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_30_5  co_30 co_i_30_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_30_6  co_30 co_i_30_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_30_7  co_30 co_i_30_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_0  co_31 co_i_31_0  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_1  co_31 co_i_31_1  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_2  co_31 co_i_31_2  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_3  co_31 co_i_31_3  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_4  co_31 co_i_31_4  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_5  co_31 co_i_31_5  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_6  co_31 co_i_31_6  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_7  co_31 co_i_31_7  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_8  co_31 co_i_31_8  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_9  co_31 co_i_31_9  VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_10 co_31 co_i_31_10 VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_11 co_31 co_i_31_11 VGND int_con C=8F R=120
x_buf1_buf16_intcon_31_12 co_31 co_i_31_12 VGND int_con C=8F R=120

x16_0_0  co_i_0_0  VGND VNB vpwr_R_1  vpwr_R_1  ff_0_0  sky130_fd_sc_hd__clkbuf_16
x16_0_1  co_i_0_1  VGND VNB vpwr_R_2  vpwr_R_2  ff_0_1  sky130_fd_sc_hd__clkbuf_16
x16_0_2  co_i_0_2  VGND VNB vpwr_R_3  vpwr_R_3  ff_0_2  sky130_fd_sc_hd__clkbuf_16
x16_0_3  co_i_0_3  VGND VNB vpwr_R_4  vpwr_R_4  ff_0_3  sky130_fd_sc_hd__clkbuf_16
x16_0_4  co_i_0_4  VGND VNB vpwr_R_5  vpwr_R_5  ff_0_4  sky130_fd_sc_hd__clkbuf_16
x16_0_5  co_i_0_5  VGND VNB vpwr_R_6  vpwr_R_6  ff_0_5  sky130_fd_sc_hd__clkbuf_16
x16_0_6  co_i_0_6  VGND VNB vpwr_R_7  vpwr_R_7  ff_0_6  sky130_fd_sc_hd__clkbuf_16
x16_0_7  co_i_0_7  VGND VNB vpwr_R_8  vpwr_R_8  ff_0_7  sky130_fd_sc_hd__clkbuf_16
x16_0_8  co_i_0_8  VGND VNB vpwr_R_9  vpwr_R_9  ff_0_8  sky130_fd_sc_hd__clkbuf_16
x16_1_0  co_i_1_0  VGND VNB vpwr_R_11 vpwr_R_11 ff_1_0  sky130_fd_sc_hd__clkbuf_16
x16_1_1  co_i_1_1  VGND VNB vpwr_R_12 vpwr_R_12 ff_1_1  sky130_fd_sc_hd__clkbuf_16
x16_1_2  co_i_1_2  VGND VNB vpwr_R_13 vpwr_R_13 ff_1_2  sky130_fd_sc_hd__clkbuf_16
x16_1_3  co_i_1_3  VGND VNB vpwr_R_14 vpwr_R_14 ff_1_3  sky130_fd_sc_hd__clkbuf_16
x16_1_4  co_i_1_4  VGND VNB vpwr_R_15 vpwr_R_15 ff_1_4  sky130_fd_sc_hd__clkbuf_16
x16_1_5  co_i_1_5  VGND VNB vpwr_R_16 vpwr_R_16 ff_1_5  sky130_fd_sc_hd__clkbuf_16
x16_1_6  co_i_1_6  VGND VNB vpwr_R_17 vpwr_R_17 ff_1_6  sky130_fd_sc_hd__clkbuf_16
x16_1_7  co_i_1_7  VGND VNB vpwr_R_18 vpwr_R_18 ff_1_7  sky130_fd_sc_hd__clkbuf_16
x16_1_8  co_i_1_8  VGND VNB vpwr_R_19 vpwr_R_19 ff_1_8  sky130_fd_sc_hd__clkbuf_16
x16_1_9  co_i_1_9  VGND VNB vpwr_R_20 vpwr_R_20 ff_1_9  sky130_fd_sc_hd__clkbuf_16
x16_1_10 co_i_1_10 VGND VNB vpwr_R_21 vpwr_R_21 ff_1_10 sky130_fd_sc_hd__clkbuf_16
x16_2_0  co_i_2_0  VGND VNB vpwr_R_23 vpwr_R_23 ff_2_0  sky130_fd_sc_hd__clkbuf_16
x16_2_1  co_i_2_1  VGND VNB vpwr_R_24 vpwr_R_24 ff_2_1  sky130_fd_sc_hd__clkbuf_16
x16_2_2  co_i_2_2  VGND VNB vpwr_R_25 vpwr_R_25 ff_2_2  sky130_fd_sc_hd__clkbuf_16
x16_2_3  co_i_2_3  VGND VNB vpwr_R_26 vpwr_R_26 ff_2_3  sky130_fd_sc_hd__clkbuf_16
x16_2_4  co_i_2_4  VGND VNB vpwr_R_27 vpwr_R_27 ff_2_4  sky130_fd_sc_hd__clkbuf_16
x16_2_5  co_i_2_5  VGND VNB vpwr_R_28 vpwr_R_28 ff_2_5  sky130_fd_sc_hd__clkbuf_16
x16_2_6  co_i_2_6  VGND VNB vpwr_R_29 vpwr_R_29 ff_2_6  sky130_fd_sc_hd__clkbuf_16
x16_2_7  co_i_2_7  VGND VNB vpwr_R_30 vpwr_R_30 ff_2_7  sky130_fd_sc_hd__clkbuf_16
x16_3_0  co_i_3_0  VGND VNB vpwr_R_32 vpwr_R_32 ff_3_0  sky130_fd_sc_hd__clkbuf_16
x16_3_1  co_i_3_1  VGND VNB vpwr_R_33 vpwr_R_33 ff_3_1  sky130_fd_sc_hd__clkbuf_16
x16_3_2  co_i_3_2  VGND VNB vpwr_R_34 vpwr_R_34 ff_3_2  sky130_fd_sc_hd__clkbuf_16
x16_3_3  co_i_3_3  VGND VNB vpwr_R_35 vpwr_R_35 ff_3_3  sky130_fd_sc_hd__clkbuf_16
x16_3_4  co_i_3_4  VGND VNB vpwr_R_36 vpwr_R_36 ff_3_4  sky130_fd_sc_hd__clkbuf_16
x16_3_5  co_i_3_5  VGND VNB vpwr_R_37 vpwr_R_37 ff_3_5  sky130_fd_sc_hd__clkbuf_16
x16_3_6  co_i_3_6  VGND VNB vpwr_R_38 vpwr_R_38 ff_3_6  sky130_fd_sc_hd__clkbuf_16
x16_3_7  co_i_3_7  VGND VNB vpwr_R_39 vpwr_R_39 ff_3_7  sky130_fd_sc_hd__clkbuf_16
x16_4_0  co_i_4_0  VGND VNB vpwr_R_41 vpwr_R_41 ff_4_0  sky130_fd_sc_hd__clkbuf_16
x16_4_1  co_i_4_1  VGND VNB vpwr_R_42 vpwr_R_42 ff_4_1  sky130_fd_sc_hd__clkbuf_16
x16_4_2  co_i_4_2  VGND VNB vpwr_R_43 vpwr_R_43 ff_4_2  sky130_fd_sc_hd__clkbuf_16
x16_4_3  co_i_4_3  VGND VNB vpwr_R_44 vpwr_R_44 ff_4_3  sky130_fd_sc_hd__clkbuf_16
x16_4_4  co_i_4_4  VGND VNB vpwr_R_45 vpwr_R_45 ff_4_4  sky130_fd_sc_hd__clkbuf_16
x16_4_5  co_i_4_5  VGND VNB vpwr_R_46 vpwr_R_46 ff_4_5  sky130_fd_sc_hd__clkbuf_16
x16_4_6  co_i_4_6  VGND VNB vpwr_R_47 vpwr_R_47 ff_4_6  sky130_fd_sc_hd__clkbuf_16
x16_4_7  co_i_4_7  VGND VNB vpwr_R_48 vpwr_R_48 ff_4_7  sky130_fd_sc_hd__clkbuf_16
x16_5_0  co_i_5_0  VGND VNB vpwr_R_50 vpwr_R_50 ff_5_0  sky130_fd_sc_hd__clkbuf_16
x16_5_1  co_i_5_1  VGND VNB vpwr_R_51 vpwr_R_51 ff_5_1  sky130_fd_sc_hd__clkbuf_16
x16_5_2  co_i_5_2  VGND VNB vpwr_R_52 vpwr_R_52 ff_5_2  sky130_fd_sc_hd__clkbuf_16
x16_5_3  co_i_5_3  VGND VNB vpwr_R_53 vpwr_R_53 ff_5_3  sky130_fd_sc_hd__clkbuf_16
x16_5_4  co_i_5_4  VGND VNB vpwr_R_54 vpwr_R_54 ff_5_4  sky130_fd_sc_hd__clkbuf_16
x16_5_5  co_i_5_5  VGND VNB vpwr_R_55 vpwr_R_55 ff_5_5  sky130_fd_sc_hd__clkbuf_16
x16_5_6  co_i_5_6  VGND VNB vpwr_R_56 vpwr_R_56 ff_5_6  sky130_fd_sc_hd__clkbuf_16
x16_5_7  co_i_5_7  VGND VNB vpwr_R_57 vpwr_R_57 ff_5_7  sky130_fd_sc_hd__clkbuf_16
x16_5_8  co_i_5_8  VGND VNB vpwr_R_58 vpwr_R_58 ff_5_8  sky130_fd_sc_hd__clkbuf_16
x16_5_9  co_i_5_9  VGND VNB vpwr_R_59 vpwr_R_59 ff_5_9  sky130_fd_sc_hd__clkbuf_16
x16_5_10 co_i_5_10 VGND VNB vpwr_R_60 vpwr_R_60 ff_5_10 sky130_fd_sc_hd__clkbuf_16
x16_5_11 co_i_5_11 VGND VNB vpwr_R_61 vpwr_R_61 ff_5_11 sky130_fd_sc_hd__clkbuf_16
x16_6_0  co_i_6_0  VGND VNB vpwr_R_63 vpwr_R_63 ff_6_0  sky130_fd_sc_hd__clkbuf_16
x16_6_1  co_i_6_1  VGND VNB vpwr_R_64 vpwr_R_64 ff_6_1  sky130_fd_sc_hd__clkbuf_16
x16_6_2  co_i_6_2  VGND VNB vpwr_R_65 vpwr_R_65 ff_6_2  sky130_fd_sc_hd__clkbuf_16
x16_6_3  co_i_6_3  VGND VNB vpwr_R_66 vpwr_R_66 ff_6_3  sky130_fd_sc_hd__clkbuf_16
x16_6_4  co_i_6_4  VGND VNB vpwr_R_67 vpwr_R_67 ff_6_4  sky130_fd_sc_hd__clkbuf_16
x16_6_5  co_i_6_5  VGND VNB vpwr_R_68 vpwr_R_68 ff_6_5  sky130_fd_sc_hd__clkbuf_16
x16_6_6  co_i_6_6  VGND VNB vpwr_R_69 vpwr_R_69 ff_6_6  sky130_fd_sc_hd__clkbuf_16
x16_6_7  co_i_6_7  VGND VNB vpwr_R_70 vpwr_R_70 ff_6_7  sky130_fd_sc_hd__clkbuf_16
x16_6_8  co_i_6_8  VGND VNB vpwr_R_71 vpwr_R_71 ff_6_8  sky130_fd_sc_hd__clkbuf_16
x16_6_9  co_i_6_9  VGND VNB vpwr_R_72 vpwr_R_72 ff_6_9  sky130_fd_sc_hd__clkbuf_16
x16_7_0  co_i_7_0  VGND VNB vpwr_R_74 vpwr_R_74 ff_7_0  sky130_fd_sc_hd__clkbuf_16
x16_7_1  co_i_7_1  VGND VNB vpwr_R_75 vpwr_R_75 ff_7_1  sky130_fd_sc_hd__clkbuf_16
x16_7_2  co_i_7_2  VGND VNB vpwr_R_76 vpwr_R_76 ff_7_2  sky130_fd_sc_hd__clkbuf_16
x16_7_3  co_i_7_3  VGND VNB vpwr_R_77 vpwr_R_77 ff_7_3  sky130_fd_sc_hd__clkbuf_16
x16_7_4  co_i_7_4  VGND VNB vpwr_R_78 vpwr_R_78 ff_7_4  sky130_fd_sc_hd__clkbuf_16
x16_7_5  co_i_7_5  VGND VNB vpwr_R_79 vpwr_R_79 ff_7_5  sky130_fd_sc_hd__clkbuf_16
x16_7_6  co_i_7_6  VGND VNB vpwr_R_80 vpwr_R_80 ff_7_6  sky130_fd_sc_hd__clkbuf_16
x16_7_7  co_i_7_7  VGND VNB vpwr_R_81 vpwr_R_81 ff_7_7  sky130_fd_sc_hd__clkbuf_16
x16_7_8  co_i_7_8  VGND VNB vpwr_R_82 vpwr_R_82 ff_7_8  sky130_fd_sc_hd__clkbuf_16
x16_7_9  co_i_7_9  VGND VNB vpwr_R_83 vpwr_R_83 ff_7_9  sky130_fd_sc_hd__clkbuf_16
x16_7_10 co_i_7_10 VGND VNB vpwr_R_84 vpwr_R_84 ff_7_10 sky130_fd_sc_hd__clkbuf_16
x16_7_11 co_i_7_11 VGND VNB vpwr_R_85 vpwr_R_85 ff_7_11 sky130_fd_sc_hd__clkbuf_16
x16_7_12 co_i_7_12 VGND VNB vpwr_R_86 vpwr_R_86 ff_7_12 sky130_fd_sc_hd__clkbuf_16
x16_7_13 co_i_7_13 VGND VNB vpwr_R_87 vpwr_R_87 ff_7_13 sky130_fd_sc_hd__clkbuf_16
x16_7_14 co_i_7_14 VGND VNB vpwr_R_88 vpwr_R_88 ff_7_14 sky130_fd_sc_hd__clkbuf_16
x16_8_0  co_i_8_0  VGND VNB vpwr_R_90 vpwr_R_90 ff_8_0  sky130_fd_sc_hd__clkbuf_16
x16_8_1  co_i_8_1  VGND VNB vpwr_R_91 vpwr_R_91 ff_8_1  sky130_fd_sc_hd__clkbuf_16
x16_8_2  co_i_8_2  VGND VNB vpwr_R_92 vpwr_R_92 ff_8_2  sky130_fd_sc_hd__clkbuf_16
x16_8_3  co_i_8_3  VGND VNB vpwr_R_93 vpwr_R_93 ff_8_3  sky130_fd_sc_hd__clkbuf_16
x16_9_0  co_i_9_0  VGND VNB vpwr_R_95 vpwr_R_95 ff_9_0  sky130_fd_sc_hd__clkbuf_16
x16_9_1  co_i_9_1  VGND VNB vpwr_R_96 vpwr_R_96 ff_9_1  sky130_fd_sc_hd__clkbuf_16
x16_9_2  co_i_9_2  VGND VNB vpwr_R_97 vpwr_R_97 ff_9_2  sky130_fd_sc_hd__clkbuf_16
x16_9_3  co_i_9_3  VGND VNB vpwr_R_98 vpwr_R_98 ff_9_3  sky130_fd_sc_hd__clkbuf_16
x16_9_4  co_i_9_4  VGND VNB vpwr_R_99 vpwr_R_99 ff_9_4  sky130_fd_sc_hd__clkbuf_16
x16_10_0  co_i_10_0  VGND VNB vpwr_R_101 vpwr_R_101 ff_10_0  sky130_fd_sc_hd__clkbuf_16
x16_10_1  co_i_10_1  VGND VNB vpwr_R_102 vpwr_R_102 ff_10_1  sky130_fd_sc_hd__clkbuf_16
x16_10_2  co_i_10_2  VGND VNB vpwr_R_103 vpwr_R_103 ff_10_2  sky130_fd_sc_hd__clkbuf_16
x16_10_3  co_i_10_3  VGND VNB vpwr_R_104 vpwr_R_104 ff_10_3  sky130_fd_sc_hd__clkbuf_16
x16_10_4  co_i_10_4  VGND VNB vpwr_R_105 vpwr_R_105 ff_10_4  sky130_fd_sc_hd__clkbuf_16
x16_10_5  co_i_10_5  VGND VNB vpwr_R_106 vpwr_R_106 ff_10_5  sky130_fd_sc_hd__clkbuf_16
x16_10_6  co_i_10_6  VGND VNB vpwr_R_107 vpwr_R_107 ff_10_6  sky130_fd_sc_hd__clkbuf_16
x16_11_0  co_i_11_0  VGND VNB vpwr_R_109 vpwr_R_109 ff_11_0  sky130_fd_sc_hd__clkbuf_16
x16_11_1  co_i_11_1  VGND VNB vpwr_R_110 vpwr_R_110 ff_11_1  sky130_fd_sc_hd__clkbuf_16
x16_11_2  co_i_11_2  VGND VNB vpwr_R_111 vpwr_R_111 ff_11_2  sky130_fd_sc_hd__clkbuf_16
x16_11_3  co_i_11_3  VGND VNB vpwr_R_112 vpwr_R_112 ff_11_3  sky130_fd_sc_hd__clkbuf_16
x16_11_4  co_i_11_4  VGND VNB vpwr_R_113 vpwr_R_113 ff_11_4  sky130_fd_sc_hd__clkbuf_16
x16_11_5  co_i_11_5  VGND VNB vpwr_R_114 vpwr_R_114 ff_11_5  sky130_fd_sc_hd__clkbuf_16
x16_11_6  co_i_11_6  VGND VNB vpwr_R_115 vpwr_R_115 ff_11_6  sky130_fd_sc_hd__clkbuf_16
x16_11_7  co_i_11_7  VGND VNB vpwr_R_116 vpwr_R_116 ff_11_7  sky130_fd_sc_hd__clkbuf_16
x16_12_0  co_i_12_0  VGND VNB vpwr_R_118 vpwr_R_118 ff_12_0  sky130_fd_sc_hd__clkbuf_16
x16_12_1  co_i_12_1  VGND VNB vpwr_R_119 vpwr_R_119 ff_12_1  sky130_fd_sc_hd__clkbuf_16
x16_12_2  co_i_12_2  VGND VNB vpwr_R_120 vpwr_R_120 ff_12_2  sky130_fd_sc_hd__clkbuf_16
x16_12_3  co_i_12_3  VGND VNB vpwr_R_121 vpwr_R_121 ff_12_3  sky130_fd_sc_hd__clkbuf_16
x16_12_4  co_i_12_4  VGND VNB vpwr_R_122 vpwr_R_122 ff_12_4  sky130_fd_sc_hd__clkbuf_16
x16_13_0  co_i_13_0  VGND VNB vpwr_R_124 vpwr_R_124 ff_13_0  sky130_fd_sc_hd__clkbuf_16
x16_13_1  co_i_13_1  VGND VNB vpwr_R_125 vpwr_R_125 ff_13_1  sky130_fd_sc_hd__clkbuf_16
x16_13_2  co_i_13_2  VGND VNB vpwr_R_126 vpwr_R_126 ff_13_2  sky130_fd_sc_hd__clkbuf_16
x16_13_3  co_i_13_3  VGND VNB vpwr_R_127 vpwr_R_127 ff_13_3  sky130_fd_sc_hd__clkbuf_16
x16_13_4  co_i_13_4  VGND VNB vpwr_R_128 vpwr_R_128 ff_13_4  sky130_fd_sc_hd__clkbuf_16
x16_13_5  co_i_13_5  VGND VNB vpwr_R_129 vpwr_R_129 ff_13_5  sky130_fd_sc_hd__clkbuf_16
x16_13_6  co_i_13_6  VGND VNB vpwr_R_130 vpwr_R_130 ff_13_6  sky130_fd_sc_hd__clkbuf_16
x16_14_0  co_i_14_0  VGND VNB vpwr_R_132 vpwr_R_132 ff_14_0  sky130_fd_sc_hd__clkbuf_16
x16_14_1  co_i_14_1  VGND VNB vpwr_R_133 vpwr_R_133 ff_14_1  sky130_fd_sc_hd__clkbuf_16
x16_14_2  co_i_14_2  VGND VNB vpwr_R_134 vpwr_R_134 ff_14_2  sky130_fd_sc_hd__clkbuf_16
x16_14_3  co_i_14_3  VGND VNB vpwr_R_135 vpwr_R_135 ff_14_3  sky130_fd_sc_hd__clkbuf_16
x16_14_4  co_i_14_4  VGND VNB vpwr_R_136 vpwr_R_136 ff_14_4  sky130_fd_sc_hd__clkbuf_16
x16_15_0  co_i_15_0  VGND VNB vpwr_R_138 vpwr_R_138 ff_15_0  sky130_fd_sc_hd__clkbuf_16
x16_15_1  co_i_15_1  VGND VNB vpwr_R_139 vpwr_R_139 ff_15_1  sky130_fd_sc_hd__clkbuf_16
x16_15_2  co_i_15_2  VGND VNB vpwr_R_140 vpwr_R_140 ff_15_2  sky130_fd_sc_hd__clkbuf_16
x16_15_3  co_i_15_3  VGND VNB vpwr_R_141 vpwr_R_141 ff_15_3  sky130_fd_sc_hd__clkbuf_16
x16_15_4  co_i_15_4  VGND VNB vpwr_R_142 vpwr_R_142 ff_15_4  sky130_fd_sc_hd__clkbuf_16
x16_15_5  co_i_15_5  VGND VNB vpwr_R_143 vpwr_R_143 ff_15_5  sky130_fd_sc_hd__clkbuf_16
x16_15_6  co_i_15_6  VGND VNB vpwr_R_144 vpwr_R_144 ff_15_6  sky130_fd_sc_hd__clkbuf_16
x16_16_0  co_i_16_0  VGND VNB vpwr_R_146 vpwr_R_146 ff_16_0  sky130_fd_sc_hd__clkbuf_16
x16_16_1  co_i_16_1  VGND VNB vpwr_R_147 vpwr_R_147 ff_16_1  sky130_fd_sc_hd__clkbuf_16
x16_16_2  co_i_16_2  VGND VNB vpwr_R_148 vpwr_R_148 ff_16_2  sky130_fd_sc_hd__clkbuf_16
x16_16_3  co_i_16_3  VGND VNB vpwr_R_149 vpwr_R_149 ff_16_3  sky130_fd_sc_hd__clkbuf_16
x16_16_4  co_i_16_4  VGND VNB vpwr_R_150 vpwr_R_150 ff_16_4  sky130_fd_sc_hd__clkbuf_16
x16_16_5  co_i_16_5  VGND VNB vpwr_R_151 vpwr_R_151 ff_16_5  sky130_fd_sc_hd__clkbuf_16
x16_16_6  co_i_16_6  VGND VNB vpwr_R_152 vpwr_R_152 ff_16_6  sky130_fd_sc_hd__clkbuf_16
x16_16_7  co_i_16_7  VGND VNB vpwr_R_153 vpwr_R_153 ff_16_7  sky130_fd_sc_hd__clkbuf_16
x16_16_8  co_i_16_8  VGND VNB vpwr_R_154 vpwr_R_154 ff_16_8  sky130_fd_sc_hd__clkbuf_16
x16_16_9  co_i_16_9  VGND VNB vpwr_R_155 vpwr_R_155 ff_16_9  sky130_fd_sc_hd__clkbuf_16
x16_16_10 co_i_16_10 VGND VNB vpwr_R_156 vpwr_R_156 ff_16_10 sky130_fd_sc_hd__clkbuf_16
x16_17_0  co_i_17_0  VGND VNB vpwr_R_158 vpwr_R_158 ff_17_0  sky130_fd_sc_hd__clkbuf_16
x16_17_1  co_i_17_1  VGND VNB vpwr_R_159 vpwr_R_159 ff_17_1  sky130_fd_sc_hd__clkbuf_16
x16_17_2  co_i_17_2  VGND VNB vpwr_R_160 vpwr_R_160 ff_17_2  sky130_fd_sc_hd__clkbuf_16
x16_17_3  co_i_17_3  VGND VNB vpwr_R_161 vpwr_R_161 ff_17_3  sky130_fd_sc_hd__clkbuf_16
x16_17_4  co_i_17_4  VGND VNB vpwr_R_162 vpwr_R_162 ff_17_4  sky130_fd_sc_hd__clkbuf_16
x16_17_5  co_i_17_5  VGND VNB vpwr_R_163 vpwr_R_163 ff_17_5  sky130_fd_sc_hd__clkbuf_16
x16_17_6  co_i_17_6  VGND VNB vpwr_R_164 vpwr_R_164 ff_17_6  sky130_fd_sc_hd__clkbuf_16
x16_17_7  co_i_17_7  VGND VNB vpwr_R_165 vpwr_R_165 ff_17_7  sky130_fd_sc_hd__clkbuf_16
x16_17_8  co_i_17_8  VGND VNB vpwr_R_166 vpwr_R_166 ff_17_8  sky130_fd_sc_hd__clkbuf_16
x16_17_9  co_i_17_9  VGND VNB vpwr_R_167 vpwr_R_167 ff_17_9  sky130_fd_sc_hd__clkbuf_16
x16_17_10 co_i_17_10 VGND VNB vpwr_R_168 vpwr_R_168 ff_17_10 sky130_fd_sc_hd__clkbuf_16
x16_17_11 co_i_17_11 VGND VNB vpwr_R_169 vpwr_R_169 ff_17_11 sky130_fd_sc_hd__clkbuf_16
x16_17_12 co_i_17_12 VGND VNB vpwr_R_170 vpwr_R_170 ff_17_12 sky130_fd_sc_hd__clkbuf_16
x16_17_13 co_i_17_13 VGND VNB vpwr_R_171 vpwr_R_171 ff_17_13 sky130_fd_sc_hd__clkbuf_16
x16_18_0  co_i_18_0  VGND VNB vpwr_R_173 vpwr_R_173 ff_18_0  sky130_fd_sc_hd__clkbuf_16
x16_18_1  co_i_18_1  VGND VNB vpwr_R_174 vpwr_R_174 ff_18_1  sky130_fd_sc_hd__clkbuf_16
x16_18_2  co_i_18_2  VGND VNB vpwr_R_175 vpwr_R_175 ff_18_2  sky130_fd_sc_hd__clkbuf_16
x16_18_3  co_i_18_3  VGND VNB vpwr_R_176 vpwr_R_176 ff_18_3  sky130_fd_sc_hd__clkbuf_16
x16_18_4  co_i_18_4  VGND VNB vpwr_R_177 vpwr_R_177 ff_18_4  sky130_fd_sc_hd__clkbuf_16
x16_18_5  co_i_18_5  VGND VNB vpwr_R_178 vpwr_R_178 ff_18_5  sky130_fd_sc_hd__clkbuf_16
x16_18_6  co_i_18_6  VGND VNB vpwr_R_179 vpwr_R_179 ff_18_6  sky130_fd_sc_hd__clkbuf_16
x16_18_7  co_i_18_7  VGND VNB vpwr_R_180 vpwr_R_180 ff_18_7  sky130_fd_sc_hd__clkbuf_16
x16_18_8  co_i_18_8  VGND VNB vpwr_R_181 vpwr_R_181 ff_18_8  sky130_fd_sc_hd__clkbuf_16
x16_18_9  co_i_18_9  VGND VNB vpwr_R_182 vpwr_R_182 ff_18_9  sky130_fd_sc_hd__clkbuf_16
x16_18_10 co_i_18_10 VGND VNB vpwr_R_183 vpwr_R_183 ff_18_10 sky130_fd_sc_hd__clkbuf_16
x16_18_11 co_i_18_11 VGND VNB vpwr_R_184 vpwr_R_184 ff_18_11 sky130_fd_sc_hd__clkbuf_16
x16_18_12 co_i_18_12 VGND VNB vpwr_R_185 vpwr_R_185 ff_18_12 sky130_fd_sc_hd__clkbuf_16
x16_19_0  co_i_19_0  VGND VNB vpwr_R_187 vpwr_R_187 ff_19_0  sky130_fd_sc_hd__clkbuf_16
x16_19_1  co_i_19_1  VGND VNB vpwr_R_188 vpwr_R_188 ff_19_1  sky130_fd_sc_hd__clkbuf_16
x16_19_2  co_i_19_2  VGND VNB vpwr_R_189 vpwr_R_189 ff_19_2  sky130_fd_sc_hd__clkbuf_16
x16_19_3  co_i_19_3  VGND VNB vpwr_R_190 vpwr_R_190 ff_19_3  sky130_fd_sc_hd__clkbuf_16
x16_19_4  co_i_19_4  VGND VNB vpwr_R_191 vpwr_R_191 ff_19_4  sky130_fd_sc_hd__clkbuf_16
x16_19_5  co_i_19_5  VGND VNB vpwr_R_192 vpwr_R_192 ff_19_5  sky130_fd_sc_hd__clkbuf_16
x16_19_6  co_i_19_6  VGND VNB vpwr_R_193 vpwr_R_193 ff_19_6  sky130_fd_sc_hd__clkbuf_16
x16_19_7  co_i_19_7  VGND VNB vpwr_R_194 vpwr_R_194 ff_19_7  sky130_fd_sc_hd__clkbuf_16
x16_20_0  co_i_20_0  VGND VNB vpwr_R_196 vpwr_R_196 ff_20_0  sky130_fd_sc_hd__clkbuf_16
x16_20_1  co_i_20_1  VGND VNB vpwr_R_197 vpwr_R_197 ff_20_1  sky130_fd_sc_hd__clkbuf_16
x16_20_2  co_i_20_2  VGND VNB vpwr_R_198 vpwr_R_198 ff_20_2  sky130_fd_sc_hd__clkbuf_16
x16_20_3  co_i_20_3  VGND VNB vpwr_R_199 vpwr_R_199 ff_20_3  sky130_fd_sc_hd__clkbuf_16
x16_20_4  co_i_20_4  VGND VNB vpwr_R_200 vpwr_R_200 ff_20_4  sky130_fd_sc_hd__clkbuf_16
x16_20_5  co_i_20_5  VGND VNB vpwr_R_201 vpwr_R_201 ff_20_5  sky130_fd_sc_hd__clkbuf_16
x16_20_6  co_i_20_6  VGND VNB vpwr_R_202 vpwr_R_202 ff_20_6  sky130_fd_sc_hd__clkbuf_16
x16_20_7  co_i_20_7  VGND VNB vpwr_R_203 vpwr_R_203 ff_20_7  sky130_fd_sc_hd__clkbuf_16
x16_20_8  co_i_20_8  VGND VNB vpwr_R_204 vpwr_R_204 ff_20_8  sky130_fd_sc_hd__clkbuf_16
x16_20_9  co_i_20_9  VGND VNB vpwr_R_205 vpwr_R_205 ff_20_9  sky130_fd_sc_hd__clkbuf_16
x16_20_10 co_i_20_10 VGND VNB vpwr_R_206 vpwr_R_206 ff_20_10 sky130_fd_sc_hd__clkbuf_16
x16_20_11 co_i_20_11 VGND VNB vpwr_R_207 vpwr_R_207 ff_20_11 sky130_fd_sc_hd__clkbuf_16
x16_20_12 co_i_20_12 VGND VNB vpwr_R_208 vpwr_R_208 ff_20_12 sky130_fd_sc_hd__clkbuf_16
x16_20_13 co_i_20_13 VGND VNB vpwr_R_209 vpwr_R_209 ff_20_13 sky130_fd_sc_hd__clkbuf_16
x16_20_14 co_i_20_14 VGND VNB vpwr_R_210 vpwr_R_210 ff_20_14 sky130_fd_sc_hd__clkbuf_16
x16_21_0  co_i_21_0  VGND VNB vpwr_R_212 vpwr_R_212 ff_21_0  sky130_fd_sc_hd__clkbuf_16
x16_21_1  co_i_21_1  VGND VNB vpwr_R_213 vpwr_R_213 ff_21_1  sky130_fd_sc_hd__clkbuf_16
x16_21_2  co_i_21_2  VGND VNB vpwr_R_214 vpwr_R_214 ff_21_2  sky130_fd_sc_hd__clkbuf_16
x16_21_3  co_i_21_3  VGND VNB vpwr_R_215 vpwr_R_215 ff_21_3  sky130_fd_sc_hd__clkbuf_16
x16_21_4  co_i_21_4  VGND VNB vpwr_R_216 vpwr_R_216 ff_21_4  sky130_fd_sc_hd__clkbuf_16
x16_21_5  co_i_21_5  VGND VNB vpwr_R_217 vpwr_R_217 ff_21_5  sky130_fd_sc_hd__clkbuf_16
x16_21_6  co_i_21_6  VGND VNB vpwr_R_218 vpwr_R_218 ff_21_6  sky130_fd_sc_hd__clkbuf_16
x16_21_7  co_i_21_7  VGND VNB vpwr_R_219 vpwr_R_219 ff_21_7  sky130_fd_sc_hd__clkbuf_16
x16_21_8  co_i_21_8  VGND VNB vpwr_R_220 vpwr_R_220 ff_21_8  sky130_fd_sc_hd__clkbuf_16
x16_21_9  co_i_21_9  VGND VNB vpwr_R_221 vpwr_R_221 ff_21_9  sky130_fd_sc_hd__clkbuf_16
x16_21_10 co_i_21_10 VGND VNB vpwr_R_222 vpwr_R_222 ff_21_10 sky130_fd_sc_hd__clkbuf_16
x16_21_11 co_i_21_11 VGND VNB vpwr_R_223 vpwr_R_223 ff_21_11 sky130_fd_sc_hd__clkbuf_16
x16_21_12 co_i_21_12 VGND VNB vpwr_R_224 vpwr_R_224 ff_21_12 sky130_fd_sc_hd__clkbuf_16
x16_22_0  co_i_22_0  VGND VNB vpwr_R_226 vpwr_R_226 ff_22_0  sky130_fd_sc_hd__clkbuf_16
x16_22_1  co_i_22_1  VGND VNB vpwr_R_227 vpwr_R_227 ff_22_1  sky130_fd_sc_hd__clkbuf_16
x16_22_2  co_i_22_2  VGND VNB vpwr_R_228 vpwr_R_228 ff_22_2  sky130_fd_sc_hd__clkbuf_16
x16_22_3  co_i_22_3  VGND VNB vpwr_R_229 vpwr_R_229 ff_22_3  sky130_fd_sc_hd__clkbuf_16
x16_22_4  co_i_22_4  VGND VNB vpwr_R_230 vpwr_R_230 ff_22_4  sky130_fd_sc_hd__clkbuf_16
x16_22_5  co_i_22_5  VGND VNB vpwr_R_231 vpwr_R_231 ff_22_5  sky130_fd_sc_hd__clkbuf_16
x16_22_6  co_i_22_6  VGND VNB vpwr_R_232 vpwr_R_232 ff_22_6  sky130_fd_sc_hd__clkbuf_16
x16_22_7  co_i_22_7  VGND VNB vpwr_R_233 vpwr_R_233 ff_22_7  sky130_fd_sc_hd__clkbuf_16
x16_22_8  co_i_22_8  VGND VNB vpwr_R_234 vpwr_R_234 ff_22_8  sky130_fd_sc_hd__clkbuf_16
x16_22_9  co_i_22_9  VGND VNB vpwr_R_235 vpwr_R_235 ff_22_9  sky130_fd_sc_hd__clkbuf_16
x16_23_0  co_i_23_0  VGND VNB vpwr_R_237 vpwr_R_237 ff_23_0  sky130_fd_sc_hd__clkbuf_16
x16_23_1  co_i_23_1  VGND VNB vpwr_R_238 vpwr_R_238 ff_23_1  sky130_fd_sc_hd__clkbuf_16
x16_23_2  co_i_23_2  VGND VNB vpwr_R_239 vpwr_R_239 ff_23_2  sky130_fd_sc_hd__clkbuf_16
x16_23_3  co_i_23_3  VGND VNB vpwr_R_240 vpwr_R_240 ff_23_3  sky130_fd_sc_hd__clkbuf_16
x16_23_4  co_i_23_4  VGND VNB vpwr_R_241 vpwr_R_241 ff_23_4  sky130_fd_sc_hd__clkbuf_16
x16_23_5  co_i_23_5  VGND VNB vpwr_R_242 vpwr_R_242 ff_23_5  sky130_fd_sc_hd__clkbuf_16
x16_23_6  co_i_23_6  VGND VNB vpwr_R_243 vpwr_R_243 ff_23_6  sky130_fd_sc_hd__clkbuf_16
x16_23_7  co_i_23_7  VGND VNB vpwr_R_244 vpwr_R_244 ff_23_7  sky130_fd_sc_hd__clkbuf_16
x16_23_8  co_i_23_8  VGND VNB vpwr_R_245 vpwr_R_245 ff_23_8  sky130_fd_sc_hd__clkbuf_16
x16_23_9  co_i_23_9  VGND VNB vpwr_R_246 vpwr_R_246 ff_23_9  sky130_fd_sc_hd__clkbuf_16
x16_23_10 co_i_23_10 VGND VNB vpwr_R_247 vpwr_R_247 ff_23_10 sky130_fd_sc_hd__clkbuf_16
x16_23_11 co_i_23_11 VGND VNB vpwr_R_248 vpwr_R_248 ff_23_11 sky130_fd_sc_hd__clkbuf_16
x16_23_12 co_i_23_12 VGND VNB vpwr_R_249 vpwr_R_249 ff_23_12 sky130_fd_sc_hd__clkbuf_16
x16_23_13 co_i_23_13 VGND VNB vpwr_R_250 vpwr_R_250 ff_23_13 sky130_fd_sc_hd__clkbuf_16
x16_23_14 co_i_23_14 VGND VNB vpwr_R_251 vpwr_R_251 ff_23_14 sky130_fd_sc_hd__clkbuf_16
x16_23_15 co_i_23_15 VGND VNB vpwr_R_252 vpwr_R_252 ff_23_15 sky130_fd_sc_hd__clkbuf_16
x16_24_0  co_i_24_0  VGND VNB vpwr_R_254 vpwr_R_254 ff_24_0  sky130_fd_sc_hd__clkbuf_16
x16_24_1  co_i_24_1  VGND VNB vpwr_R_255 vpwr_R_255 ff_24_1  sky130_fd_sc_hd__clkbuf_16
x16_24_2  co_i_24_2  VGND VNB vpwr_R_256 vpwr_R_256 ff_24_2  sky130_fd_sc_hd__clkbuf_16
x16_24_3  co_i_24_3  VGND VNB vpwr_R_257 vpwr_R_257 ff_24_3  sky130_fd_sc_hd__clkbuf_16
x16_24_4  co_i_24_4  VGND VNB vpwr_R_258 vpwr_R_258 ff_24_4  sky130_fd_sc_hd__clkbuf_16
x16_24_5  co_i_24_5  VGND VNB vpwr_R_259 vpwr_R_259 ff_24_5  sky130_fd_sc_hd__clkbuf_16
x16_24_6  co_i_24_6  VGND VNB vpwr_R_260 vpwr_R_260 ff_24_6  sky130_fd_sc_hd__clkbuf_16
x16_24_7  co_i_24_7  VGND VNB vpwr_R_261 vpwr_R_261 ff_24_7  sky130_fd_sc_hd__clkbuf_16
x16_24_8  co_i_24_8  VGND VNB vpwr_R_262 vpwr_R_262 ff_24_8  sky130_fd_sc_hd__clkbuf_16
x16_24_9  co_i_24_9  VGND VNB vpwr_R_263 vpwr_R_263 ff_24_9  sky130_fd_sc_hd__clkbuf_16
x16_24_10 co_i_24_10 VGND VNB vpwr_R_264 vpwr_R_264 ff_24_10 sky130_fd_sc_hd__clkbuf_16
x16_25_0  co_i_25_0  VGND VNB vpwr_R_266 vpwr_R_266 ff_25_0  sky130_fd_sc_hd__clkbuf_16
x16_25_1  co_i_25_1  VGND VNB vpwr_R_267 vpwr_R_267 ff_25_1  sky130_fd_sc_hd__clkbuf_16
x16_25_2  co_i_25_2  VGND VNB vpwr_R_268 vpwr_R_268 ff_25_2  sky130_fd_sc_hd__clkbuf_16
x16_25_3  co_i_25_3  VGND VNB vpwr_R_269 vpwr_R_269 ff_25_3  sky130_fd_sc_hd__clkbuf_16
x16_25_4  co_i_25_4  VGND VNB vpwr_R_270 vpwr_R_270 ff_25_4  sky130_fd_sc_hd__clkbuf_16
x16_25_5  co_i_25_5  VGND VNB vpwr_R_271 vpwr_R_271 ff_25_5  sky130_fd_sc_hd__clkbuf_16
x16_25_6  co_i_25_6  VGND VNB vpwr_R_272 vpwr_R_272 ff_25_6  sky130_fd_sc_hd__clkbuf_16
x16_25_7  co_i_25_7  VGND VNB vpwr_R_273 vpwr_R_273 ff_25_7  sky130_fd_sc_hd__clkbuf_16
x16_25_8  co_i_25_8  VGND VNB vpwr_R_274 vpwr_R_274 ff_25_8  sky130_fd_sc_hd__clkbuf_16
x16_25_9  co_i_25_9  VGND VNB vpwr_R_275 vpwr_R_275 ff_25_9  sky130_fd_sc_hd__clkbuf_16
x16_25_10 co_i_25_10 VGND VNB vpwr_R_276 vpwr_R_276 ff_25_10 sky130_fd_sc_hd__clkbuf_16
x16_25_11 co_i_25_11 VGND VNB vpwr_R_277 vpwr_R_277 ff_25_11 sky130_fd_sc_hd__clkbuf_16
x16_26_0  co_i_26_0  VGND VNB vpwr_R_279 vpwr_R_279 ff_26_0  sky130_fd_sc_hd__clkbuf_16
x16_26_1  co_i_26_1  VGND VNB vpwr_R_280 vpwr_R_280 ff_26_1  sky130_fd_sc_hd__clkbuf_16
x16_26_2  co_i_26_2  VGND VNB vpwr_R_281 vpwr_R_281 ff_26_2  sky130_fd_sc_hd__clkbuf_16
x16_26_3  co_i_26_3  VGND VNB vpwr_R_282 vpwr_R_282 ff_26_3  sky130_fd_sc_hd__clkbuf_16
x16_26_4  co_i_26_4  VGND VNB vpwr_R_283 vpwr_R_283 ff_26_4  sky130_fd_sc_hd__clkbuf_16
x16_26_5  co_i_26_5  VGND VNB vpwr_R_284 vpwr_R_284 ff_26_5  sky130_fd_sc_hd__clkbuf_16
x16_26_6  co_i_26_6  VGND VNB vpwr_R_285 vpwr_R_285 ff_26_6  sky130_fd_sc_hd__clkbuf_16
x16_26_7  co_i_26_7  VGND VNB vpwr_R_286 vpwr_R_286 ff_26_7  sky130_fd_sc_hd__clkbuf_16
x16_26_8  co_i_26_8  VGND VNB vpwr_R_287 vpwr_R_287 ff_26_8  sky130_fd_sc_hd__clkbuf_16
x16_26_9  co_i_26_9  VGND VNB vpwr_R_288 vpwr_R_288 ff_26_9  sky130_fd_sc_hd__clkbuf_16
x16_27_0  co_i_27_0  VGND VNB vpwr_R_290 vpwr_R_290 ff_27_0  sky130_fd_sc_hd__clkbuf_16
x16_27_1  co_i_27_1  VGND VNB vpwr_R_291 vpwr_R_291 ff_27_1  sky130_fd_sc_hd__clkbuf_16
x16_27_2  co_i_27_2  VGND VNB vpwr_R_292 vpwr_R_292 ff_27_2  sky130_fd_sc_hd__clkbuf_16
x16_27_3  co_i_27_3  VGND VNB vpwr_R_293 vpwr_R_293 ff_27_3  sky130_fd_sc_hd__clkbuf_16
x16_27_4  co_i_27_4  VGND VNB vpwr_R_294 vpwr_R_294 ff_27_4  sky130_fd_sc_hd__clkbuf_16
x16_27_5  co_i_27_5  VGND VNB vpwr_R_295 vpwr_R_295 ff_27_5  sky130_fd_sc_hd__clkbuf_16
x16_27_6  co_i_27_6  VGND VNB vpwr_R_296 vpwr_R_296 ff_27_6  sky130_fd_sc_hd__clkbuf_16
x16_27_7  co_i_27_7  VGND VNB vpwr_R_297 vpwr_R_297 ff_27_7  sky130_fd_sc_hd__clkbuf_16
x16_27_8  co_i_27_8  VGND VNB vpwr_R_298 vpwr_R_298 ff_27_8  sky130_fd_sc_hd__clkbuf_16
x16_28_0  co_i_28_0  VGND VNB vpwr_R_300 vpwr_R_300 ff_28_0  sky130_fd_sc_hd__clkbuf_16
x16_28_1  co_i_28_1  VGND VNB vpwr_R_301 vpwr_R_301 ff_28_1  sky130_fd_sc_hd__clkbuf_16
x16_28_2  co_i_28_2  VGND VNB vpwr_R_302 vpwr_R_302 ff_28_2  sky130_fd_sc_hd__clkbuf_16
x16_28_3  co_i_28_3  VGND VNB vpwr_R_303 vpwr_R_303 ff_28_3  sky130_fd_sc_hd__clkbuf_16
x16_28_4  co_i_28_4  VGND VNB vpwr_R_304 vpwr_R_304 ff_28_4  sky130_fd_sc_hd__clkbuf_16
x16_28_5  co_i_28_5  VGND VNB vpwr_R_305 vpwr_R_305 ff_28_5  sky130_fd_sc_hd__clkbuf_16
x16_28_6  co_i_28_6  VGND VNB vpwr_R_306 vpwr_R_306 ff_28_6  sky130_fd_sc_hd__clkbuf_16
x16_28_7  co_i_28_7  VGND VNB vpwr_R_307 vpwr_R_307 ff_28_7  sky130_fd_sc_hd__clkbuf_16
x16_28_8  co_i_28_8  VGND VNB vpwr_R_308 vpwr_R_308 ff_28_8  sky130_fd_sc_hd__clkbuf_16
x16_28_9  co_i_28_9  VGND VNB vpwr_R_309 vpwr_R_309 ff_28_9  sky130_fd_sc_hd__clkbuf_16
x16_28_10 co_i_28_10 VGND VNB vpwr_R_310 vpwr_R_310 ff_28_10 sky130_fd_sc_hd__clkbuf_16
x16_28_11 co_i_28_11 VGND VNB vpwr_R_311 vpwr_R_311 ff_28_11 sky130_fd_sc_hd__clkbuf_16
x16_28_12 co_i_28_12 VGND VNB vpwr_R_312 vpwr_R_312 ff_28_12 sky130_fd_sc_hd__clkbuf_16
x16_29_0  co_i_29_0  VGND VNB vpwr_R_314 vpwr_R_314 ff_29_0  sky130_fd_sc_hd__clkbuf_16
x16_29_1  co_i_29_1  VGND VNB vpwr_R_315 vpwr_R_315 ff_29_1  sky130_fd_sc_hd__clkbuf_16
x16_29_2  co_i_29_2  VGND VNB vpwr_R_316 vpwr_R_316 ff_29_2  sky130_fd_sc_hd__clkbuf_16
x16_29_3  co_i_29_3  VGND VNB vpwr_R_317 vpwr_R_317 ff_29_3  sky130_fd_sc_hd__clkbuf_16
x16_29_4  co_i_29_4  VGND VNB vpwr_R_318 vpwr_R_318 ff_29_4  sky130_fd_sc_hd__clkbuf_16
x16_29_5  co_i_29_5  VGND VNB vpwr_R_319 vpwr_R_319 ff_29_5  sky130_fd_sc_hd__clkbuf_16
x16_29_6  co_i_29_6  VGND VNB vpwr_R_320 vpwr_R_320 ff_29_6  sky130_fd_sc_hd__clkbuf_16
x16_29_7  co_i_29_7  VGND VNB vpwr_R_321 vpwr_R_321 ff_29_7  sky130_fd_sc_hd__clkbuf_16
x16_29_8  co_i_29_8  VGND VNB vpwr_R_322 vpwr_R_322 ff_29_8  sky130_fd_sc_hd__clkbuf_16
x16_29_9  co_i_29_9  VGND VNB vpwr_R_323 vpwr_R_323 ff_29_9  sky130_fd_sc_hd__clkbuf_16
x16_29_10 co_i_29_10 VGND VNB vpwr_R_324 vpwr_R_324 ff_29_10 sky130_fd_sc_hd__clkbuf_16
x16_29_11 co_i_29_11 VGND VNB vpwr_R_325 vpwr_R_325 ff_29_11 sky130_fd_sc_hd__clkbuf_16
x16_29_12 co_i_29_12 VGND VNB vpwr_R_326 vpwr_R_326 ff_29_12 sky130_fd_sc_hd__clkbuf_16
x16_30_0  co_i_30_0  VGND VNB vpwr_R_328 vpwr_R_328 ff_30_0  sky130_fd_sc_hd__clkbuf_16
x16_30_1  co_i_30_1  VGND VNB vpwr_R_329 vpwr_R_329 ff_30_1  sky130_fd_sc_hd__clkbuf_16
x16_30_2  co_i_30_2  VGND VNB vpwr_R_330 vpwr_R_330 ff_30_2  sky130_fd_sc_hd__clkbuf_16
x16_30_3  co_i_30_3  VGND VNB vpwr_R_331 vpwr_R_331 ff_30_3  sky130_fd_sc_hd__clkbuf_16
x16_30_4  co_i_30_4  VGND VNB vpwr_R_332 vpwr_R_332 ff_30_4  sky130_fd_sc_hd__clkbuf_16
x16_30_5  co_i_30_5  VGND VNB vpwr_R_333 vpwr_R_333 ff_30_5  sky130_fd_sc_hd__clkbuf_16
x16_30_6  co_i_30_6  VGND VNB vpwr_R_334 vpwr_R_334 ff_30_6  sky130_fd_sc_hd__clkbuf_16
x16_30_7  co_i_30_7  VGND VNB vpwr_R_335 vpwr_R_335 ff_30_7  sky130_fd_sc_hd__clkbuf_16
x16_31_0  co_i_31_0  VGND VNB vpwr_R_337 vpwr_R_337 ff_31_0  sky130_fd_sc_hd__clkbuf_16
x16_31_1  co_i_31_1  VGND VNB vpwr_R_338 vpwr_R_338 ff_31_1  sky130_fd_sc_hd__clkbuf_16
x16_31_2  co_i_31_2  VGND VNB vpwr_R_339 vpwr_R_339 ff_31_2  sky130_fd_sc_hd__clkbuf_16
x16_31_3  co_i_31_3  VGND VNB vpwr_R_340 vpwr_R_340 ff_31_3  sky130_fd_sc_hd__clkbuf_16
x16_31_4  co_i_31_4  VGND VNB vpwr_R_341 vpwr_R_341 ff_31_4  sky130_fd_sc_hd__clkbuf_16
x16_31_5  co_i_31_5  VGND VNB vpwr_R_342 vpwr_R_342 ff_31_5  sky130_fd_sc_hd__clkbuf_16
x16_31_6  co_i_31_6  VGND VNB vpwr_R_343 vpwr_R_343 ff_31_6  sky130_fd_sc_hd__clkbuf_16
x16_31_7  co_i_31_7  VGND VNB vpwr_R_344 vpwr_R_344 ff_31_7  sky130_fd_sc_hd__clkbuf_16
x16_31_8  co_i_31_8  VGND VNB vpwr_R_345 vpwr_R_345 ff_31_8  sky130_fd_sc_hd__clkbuf_16
x16_31_9  co_i_31_9  VGND VNB vpwr_R_346 vpwr_R_346 ff_31_9  sky130_fd_sc_hd__clkbuf_16
x16_31_10 co_i_31_10 VGND VNB vpwr_R_347 vpwr_R_347 ff_31_10 sky130_fd_sc_hd__clkbuf_16
x16_31_11 co_i_31_11 VGND VNB vpwr_R_348 vpwr_R_348 ff_31_11 sky130_fd_sc_hd__clkbuf_16
x16_31_12 co_i_31_12 VGND VNB vpwr_R_349 vpwr_R_349 ff_31_12 sky130_fd_sc_hd__clkbuf_16

xf_0_0  ff_0_0  ff_clk_0_0  VGND ff_rc m=11
xf_0_1  ff_0_1  ff_clk_0_1  VGND ff_rc m=15
xf_0_2  ff_0_2  ff_clk_0_2  VGND ff_rc m=10
xf_0_3  ff_0_3  ff_clk_0_3  VGND ff_rc m=14
xf_0_4  ff_0_4  ff_clk_0_4  VGND ff_rc m=9
xf_0_5  ff_0_5  ff_clk_0_5  VGND ff_rc m=10
xf_0_6  ff_0_6  ff_clk_0_6  VGND ff_rc m=5
xf_0_7  ff_0_7  ff_clk_0_7  VGND ff_rc m=15
xf_0_8  ff_0_8  ff_clk_0_8  VGND ff_rc m=9
xf_1_0  ff_1_0  ff_clk_1_0  VGND ff_rc m=14
xf_1_1  ff_1_1  ff_clk_1_1  VGND ff_rc m=8
xf_1_2  ff_1_2  ff_clk_1_2  VGND ff_rc m=15
xf_1_3  ff_1_3  ff_clk_1_3  VGND ff_rc m=15
xf_1_4  ff_1_4  ff_clk_1_4  VGND ff_rc m=14
xf_1_5  ff_1_5  ff_clk_1_5  VGND ff_rc m=8
xf_1_6  ff_1_6  ff_clk_1_6  VGND ff_rc m=11
xf_1_7  ff_1_7  ff_clk_1_7  VGND ff_rc m=8
xf_1_8  ff_1_8  ff_clk_1_8  VGND ff_rc m=12
xf_1_9  ff_1_9  ff_clk_1_9  VGND ff_rc m=13
xf_1_10 ff_1_10 ff_clk_1_10 VGND ff_rc m=17
xf_2_0  ff_2_0  ff_clk_2_0  VGND ff_rc m=8
xf_2_1  ff_2_1  ff_clk_2_1  VGND ff_rc m=13
xf_2_2  ff_2_2  ff_clk_2_2  VGND ff_rc m=15
xf_2_3  ff_2_3  ff_clk_2_3  VGND ff_rc m=13
xf_2_4  ff_2_4  ff_clk_2_4  VGND ff_rc m=3
xf_2_5  ff_2_5  ff_clk_2_5  VGND ff_rc m=15
xf_2_6  ff_2_6  ff_clk_2_6  VGND ff_rc m=17
xf_2_7  ff_2_7  ff_clk_2_7  VGND ff_rc m=9
xf_3_0  ff_3_0  ff_clk_3_0  VGND ff_rc m=6
xf_3_1  ff_3_1  ff_clk_3_1  VGND ff_rc m=16
xf_3_2  ff_3_2  ff_clk_3_2  VGND ff_rc m=14
xf_3_3  ff_3_3  ff_clk_3_3  VGND ff_rc m=8
xf_3_4  ff_3_4  ff_clk_3_4  VGND ff_rc m=12
xf_3_5  ff_3_5  ff_clk_3_5  VGND ff_rc m=15
xf_3_6  ff_3_6  ff_clk_3_6  VGND ff_rc m=6
xf_3_7  ff_3_7  ff_clk_3_7  VGND ff_rc m=17
xf_4_0  ff_4_0  ff_clk_4_0  VGND ff_rc m=5
xf_4_1  ff_4_1  ff_clk_4_1  VGND ff_rc m=13
xf_4_2  ff_4_2  ff_clk_4_2  VGND ff_rc m=6
xf_4_3  ff_4_3  ff_clk_4_3  VGND ff_rc m=5
xf_4_4  ff_4_4  ff_clk_4_4  VGND ff_rc m=13
xf_4_5  ff_4_5  ff_clk_4_5  VGND ff_rc m=9
xf_4_6  ff_4_6  ff_clk_4_6  VGND ff_rc m=11
xf_4_7  ff_4_7  ff_clk_4_7  VGND ff_rc m=13
xf_5_0  ff_5_0  ff_clk_5_0  VGND ff_rc m=13
xf_5_1  ff_5_1  ff_clk_5_1  VGND ff_rc m=19
xf_5_2  ff_5_2  ff_clk_5_2  VGND ff_rc m=20
xf_5_3  ff_5_3  ff_clk_5_3  VGND ff_rc m=11
xf_5_4  ff_5_4  ff_clk_5_4  VGND ff_rc m=9
xf_5_5  ff_5_5  ff_clk_5_5  VGND ff_rc m=15
xf_5_6  ff_5_6  ff_clk_5_6  VGND ff_rc m=14
xf_5_7  ff_5_7  ff_clk_5_7  VGND ff_rc m=12
xf_5_8  ff_5_8  ff_clk_5_8  VGND ff_rc m=5
xf_5_9  ff_5_9  ff_clk_5_9  VGND ff_rc m=12
xf_5_10 ff_5_10 ff_clk_5_10 VGND ff_rc m=9
xf_5_11 ff_5_11 ff_clk_5_11 VGND ff_rc m=13
xf_6_0  ff_6_0  ff_clk_6_0  VGND ff_rc m=6
xf_6_1  ff_6_1  ff_clk_6_1  VGND ff_rc m=8
xf_6_2  ff_6_2  ff_clk_6_2  VGND ff_rc m=11
xf_6_3  ff_6_3  ff_clk_6_3  VGND ff_rc m=6
xf_6_4  ff_6_4  ff_clk_6_4  VGND ff_rc m=9
xf_6_5  ff_6_5  ff_clk_6_5  VGND ff_rc m=19
xf_6_6  ff_6_6  ff_clk_6_6  VGND ff_rc m=9
xf_6_7  ff_6_7  ff_clk_6_7  VGND ff_rc m=9
xf_6_8  ff_6_8  ff_clk_6_8  VGND ff_rc m=12
xf_6_9  ff_6_9  ff_clk_6_9  VGND ff_rc m=10
xf_7_0  ff_7_0  ff_clk_7_0  VGND ff_rc m=17
xf_7_1  ff_7_1  ff_clk_7_1  VGND ff_rc m=16
xf_7_2  ff_7_2  ff_clk_7_2  VGND ff_rc m=9
xf_7_3  ff_7_3  ff_clk_7_3  VGND ff_rc m=17
xf_7_4  ff_7_4  ff_clk_7_4  VGND ff_rc m=8
xf_7_5  ff_7_5  ff_clk_7_5  VGND ff_rc m=14
xf_7_6  ff_7_6  ff_clk_7_6  VGND ff_rc m=11
xf_7_7  ff_7_7  ff_clk_7_7  VGND ff_rc m=12
xf_7_8  ff_7_8  ff_clk_7_8  VGND ff_rc m=12
xf_7_9  ff_7_9  ff_clk_7_9  VGND ff_rc m=12
xf_7_10 ff_7_10 ff_clk_7_10 VGND ff_rc m=11
xf_7_11 ff_7_11 ff_clk_7_11 VGND ff_rc m=11
xf_7_12 ff_7_12 ff_clk_7_12 VGND ff_rc m=8
xf_7_13 ff_7_13 ff_clk_7_13 VGND ff_rc m=9
xf_7_14 ff_7_14 ff_clk_7_14 VGND ff_rc m=18
xf_8_0  ff_8_0  ff_clk_8_0  VGND ff_rc m=9
xf_8_1  ff_8_1  ff_clk_8_1  VGND ff_rc m=8
xf_8_2  ff_8_2  ff_clk_8_2  VGND ff_rc m=15
xf_8_3  ff_8_3  ff_clk_8_3  VGND ff_rc m=4
xf_9_0  ff_9_0  ff_clk_9_0  VGND ff_rc m=10
xf_9_1  ff_9_1  ff_clk_9_1  VGND ff_rc m=8
xf_9_2  ff_9_2  ff_clk_9_2  VGND ff_rc m=4
xf_9_3  ff_9_3  ff_clk_9_3  VGND ff_rc m=14
xf_9_4  ff_9_4  ff_clk_9_4  VGND ff_rc m=7
xf_10_0  ff_10_0  ff_clk_10_0  VGND ff_rc m=3
xf_10_1  ff_10_1  ff_clk_10_1  VGND ff_rc m=3
xf_10_2  ff_10_2  ff_clk_10_2  VGND ff_rc m=6
xf_10_3  ff_10_3  ff_clk_10_3  VGND ff_rc m=2
xf_10_4  ff_10_4  ff_clk_10_4  VGND ff_rc m=8
xf_10_5  ff_10_5  ff_clk_10_5  VGND ff_rc m=13
xf_10_6  ff_10_6  ff_clk_10_6  VGND ff_rc m=4
xf_11_0  ff_11_0  ff_clk_11_0  VGND ff_rc m=5
xf_11_1  ff_11_1  ff_clk_11_1  VGND ff_rc m=13
xf_11_2  ff_11_2  ff_clk_11_2  VGND ff_rc m=16
xf_11_3  ff_11_3  ff_clk_11_3  VGND ff_rc m=16
xf_11_4  ff_11_4  ff_clk_11_4  VGND ff_rc m=5
xf_11_5  ff_11_5  ff_clk_11_5  VGND ff_rc m=7
xf_11_6  ff_11_6  ff_clk_11_6  VGND ff_rc m=11
xf_11_7  ff_11_7  ff_clk_11_7  VGND ff_rc m=11
xf_12_0  ff_12_0  ff_clk_12_0  VGND ff_rc m=14
xf_12_1  ff_12_1  ff_clk_12_1  VGND ff_rc m=20
xf_12_2  ff_12_2  ff_clk_12_2  VGND ff_rc m=7
xf_12_3  ff_12_3  ff_clk_12_3  VGND ff_rc m=12
xf_12_4  ff_12_4  ff_clk_12_4  VGND ff_rc m=10
xf_13_0  ff_13_0  ff_clk_13_0  VGND ff_rc m=9
xf_13_1  ff_13_1  ff_clk_13_1  VGND ff_rc m=6
xf_13_2  ff_13_2  ff_clk_13_2  VGND ff_rc m=7
xf_13_3  ff_13_3  ff_clk_13_3  VGND ff_rc m=8
xf_13_4  ff_13_4  ff_clk_13_4  VGND ff_rc m=8
xf_13_5  ff_13_5  ff_clk_13_5  VGND ff_rc m=15
xf_13_6  ff_13_6  ff_clk_13_6  VGND ff_rc m=10
xf_14_0  ff_14_0  ff_clk_14_0  VGND ff_rc m=15
xf_14_1  ff_14_1  ff_clk_14_1  VGND ff_rc m=11
xf_14_2  ff_14_2  ff_clk_14_2  VGND ff_rc m=5
xf_14_3  ff_14_3  ff_clk_14_3  VGND ff_rc m=15
xf_14_4  ff_14_4  ff_clk_14_4  VGND ff_rc m=2
xf_15_0  ff_15_0  ff_clk_15_0  VGND ff_rc m=5
xf_15_1  ff_15_1  ff_clk_15_1  VGND ff_rc m=4
xf_15_2  ff_15_2  ff_clk_15_2  VGND ff_rc m=10
xf_15_3  ff_15_3  ff_clk_15_3  VGND ff_rc m=7
xf_15_4  ff_15_4  ff_clk_15_4  VGND ff_rc m=12
xf_15_5  ff_15_5  ff_clk_15_5  VGND ff_rc m=14
xf_15_6  ff_15_6  ff_clk_15_6  VGND ff_rc m=16
xf_16_0  ff_16_0  ff_clk_16_0  VGND ff_rc m=15
xf_16_1  ff_16_1  ff_clk_16_1  VGND ff_rc m=10
xf_16_2  ff_16_2  ff_clk_16_2  VGND ff_rc m=5
xf_16_3  ff_16_3  ff_clk_16_3  VGND ff_rc m=4
xf_16_4  ff_16_4  ff_clk_16_4  VGND ff_rc m=11
xf_16_5  ff_16_5  ff_clk_16_5  VGND ff_rc m=15
xf_16_6  ff_16_6  ff_clk_16_6  VGND ff_rc m=8
xf_16_7  ff_16_7  ff_clk_16_7  VGND ff_rc m=16
xf_16_8  ff_16_8  ff_clk_16_8  VGND ff_rc m=12
xf_16_9  ff_16_9  ff_clk_16_9  VGND ff_rc m=16
xf_16_10 ff_16_10 ff_clk_16_10 VGND ff_rc m=6
xf_17_0  ff_17_0  ff_clk_17_0  VGND ff_rc m=12
xf_17_1  ff_17_1  ff_clk_17_1  VGND ff_rc m=17
xf_17_2  ff_17_2  ff_clk_17_2  VGND ff_rc m=17
xf_17_3  ff_17_3  ff_clk_17_3  VGND ff_rc m=15
xf_17_4  ff_17_4  ff_clk_17_4  VGND ff_rc m=17
xf_17_5  ff_17_5  ff_clk_17_5  VGND ff_rc m=13
xf_17_6  ff_17_6  ff_clk_17_6  VGND ff_rc m=9
xf_17_7  ff_17_7  ff_clk_17_7  VGND ff_rc m=8
xf_17_8  ff_17_8  ff_clk_17_8  VGND ff_rc m=11
xf_17_9  ff_17_9  ff_clk_17_9  VGND ff_rc m=8
xf_17_10 ff_17_10 ff_clk_17_10 VGND ff_rc m=14
xf_17_11 ff_17_11 ff_clk_17_11 VGND ff_rc m=8
xf_17_12 ff_17_12 ff_clk_17_12 VGND ff_rc m=17
xf_17_13 ff_17_13 ff_clk_17_13 VGND ff_rc m=3
xf_18_0  ff_18_0  ff_clk_18_0  VGND ff_rc m=5
xf_18_1  ff_18_1  ff_clk_18_1  VGND ff_rc m=8
xf_18_2  ff_18_2  ff_clk_18_2  VGND ff_rc m=12
xf_18_3  ff_18_3  ff_clk_18_3  VGND ff_rc m=20
xf_18_4  ff_18_4  ff_clk_18_4  VGND ff_rc m=11
xf_18_5  ff_18_5  ff_clk_18_5  VGND ff_rc m=4
xf_18_6  ff_18_6  ff_clk_18_6  VGND ff_rc m=10
xf_18_7  ff_18_7  ff_clk_18_7  VGND ff_rc m=12
xf_18_8  ff_18_8  ff_clk_18_8  VGND ff_rc m=11
xf_18_9  ff_18_9  ff_clk_18_9  VGND ff_rc m=16
xf_18_10 ff_18_10 ff_clk_18_10 VGND ff_rc m=15
xf_18_11 ff_18_11 ff_clk_18_11 VGND ff_rc m=5
xf_18_12 ff_18_12 ff_clk_18_12 VGND ff_rc m=6
xf_19_0  ff_19_0  ff_clk_19_0  VGND ff_rc m=10
xf_19_1  ff_19_1  ff_clk_19_1  VGND ff_rc m=8
xf_19_2  ff_19_2  ff_clk_19_2  VGND ff_rc m=4
xf_19_3  ff_19_3  ff_clk_19_3  VGND ff_rc m=9
xf_19_4  ff_19_4  ff_clk_19_4  VGND ff_rc m=10
xf_19_5  ff_19_5  ff_clk_19_5  VGND ff_rc m=7
xf_19_6  ff_19_6  ff_clk_19_6  VGND ff_rc m=14
xf_19_7  ff_19_7  ff_clk_19_7  VGND ff_rc m=9
xf_20_0  ff_20_0  ff_clk_20_0  VGND ff_rc m=11
xf_20_1  ff_20_1  ff_clk_20_1  VGND ff_rc m=7
xf_20_2  ff_20_2  ff_clk_20_2  VGND ff_rc m=16
xf_20_3  ff_20_3  ff_clk_20_3  VGND ff_rc m=12
xf_20_4  ff_20_4  ff_clk_20_4  VGND ff_rc m=11
xf_20_5  ff_20_5  ff_clk_20_5  VGND ff_rc m=7
xf_20_6  ff_20_6  ff_clk_20_6  VGND ff_rc m=19
xf_20_7  ff_20_7  ff_clk_20_7  VGND ff_rc m=10
xf_20_8  ff_20_8  ff_clk_20_8  VGND ff_rc m=5
xf_20_9  ff_20_9  ff_clk_20_9  VGND ff_rc m=14
xf_20_10 ff_20_10 ff_clk_20_10 VGND ff_rc m=9
xf_20_11 ff_20_11 ff_clk_20_11 VGND ff_rc m=17
xf_20_12 ff_20_12 ff_clk_20_12 VGND ff_rc m=9
xf_20_13 ff_20_13 ff_clk_20_13 VGND ff_rc m=11
xf_20_14 ff_20_14 ff_clk_20_14 VGND ff_rc m=8
xf_21_0  ff_21_0  ff_clk_21_0  VGND ff_rc m=19
xf_21_1  ff_21_1  ff_clk_21_1  VGND ff_rc m=12
xf_21_2  ff_21_2  ff_clk_21_2  VGND ff_rc m=12
xf_21_3  ff_21_3  ff_clk_21_3  VGND ff_rc m=13
xf_21_4  ff_21_4  ff_clk_21_4  VGND ff_rc m=12
xf_21_5  ff_21_5  ff_clk_21_5  VGND ff_rc m=15
xf_21_6  ff_21_6  ff_clk_21_6  VGND ff_rc m=12
xf_21_7  ff_21_7  ff_clk_21_7  VGND ff_rc m=17
xf_21_8  ff_21_8  ff_clk_21_8  VGND ff_rc m=14
xf_21_9  ff_21_9  ff_clk_21_9  VGND ff_rc m=12
xf_21_10 ff_21_10 ff_clk_21_10 VGND ff_rc m=10
xf_21_11 ff_21_11 ff_clk_21_11 VGND ff_rc m=11
xf_21_12 ff_21_12 ff_clk_21_12 VGND ff_rc m=13
xf_22_0  ff_22_0  ff_clk_22_0  VGND ff_rc m=10
xf_22_1  ff_22_1  ff_clk_22_1  VGND ff_rc m=11
xf_22_2  ff_22_2  ff_clk_22_2  VGND ff_rc m=5
xf_22_3  ff_22_3  ff_clk_22_3  VGND ff_rc m=6
xf_22_4  ff_22_4  ff_clk_22_4  VGND ff_rc m=11
xf_22_5  ff_22_5  ff_clk_22_5  VGND ff_rc m=16
xf_22_6  ff_22_6  ff_clk_22_6  VGND ff_rc m=7
xf_22_7  ff_22_7  ff_clk_22_7  VGND ff_rc m=6
xf_22_8  ff_22_8  ff_clk_22_8  VGND ff_rc m=2
xf_22_9  ff_22_9  ff_clk_22_9  VGND ff_rc m=14
xf_23_0  ff_23_0  ff_clk_23_0  VGND ff_rc m=9
xf_23_1  ff_23_1  ff_clk_23_1  VGND ff_rc m=12
xf_23_2  ff_23_2  ff_clk_23_2  VGND ff_rc m=12
xf_23_3  ff_23_3  ff_clk_23_3  VGND ff_rc m=12
xf_23_4  ff_23_4  ff_clk_23_4  VGND ff_rc m=18
xf_23_5  ff_23_5  ff_clk_23_5  VGND ff_rc m=12
xf_23_6  ff_23_6  ff_clk_23_6  VGND ff_rc m=12
xf_23_7  ff_23_7  ff_clk_23_7  VGND ff_rc m=15
xf_23_8  ff_23_8  ff_clk_23_8  VGND ff_rc m=8
xf_23_9  ff_23_9  ff_clk_23_9  VGND ff_rc m=8
xf_23_10 ff_23_10 ff_clk_23_10 VGND ff_rc m=19
xf_23_11 ff_23_11 ff_clk_23_11 VGND ff_rc m=7
xf_23_12 ff_23_12 ff_clk_23_12 VGND ff_rc m=6
xf_23_13 ff_23_13 ff_clk_23_13 VGND ff_rc m=10
xf_23_14 ff_23_14 ff_clk_23_14 VGND ff_rc m=9
xf_23_15 ff_23_15 ff_clk_23_15 VGND ff_rc m=10
xf_24_0  ff_24_0  ff_clk_24_0  VGND ff_rc m=8
xf_24_1  ff_24_1  ff_clk_24_1  VGND ff_rc m=17
xf_24_2  ff_24_2  ff_clk_24_2  VGND ff_rc m=14
xf_24_3  ff_24_3  ff_clk_24_3  VGND ff_rc m=18
xf_24_4  ff_24_4  ff_clk_24_4  VGND ff_rc m=9
xf_24_5  ff_24_5  ff_clk_24_5  VGND ff_rc m=7
xf_24_6  ff_24_6  ff_clk_24_6  VGND ff_rc m=14
xf_24_7  ff_24_7  ff_clk_24_7  VGND ff_rc m=20
xf_24_8  ff_24_8  ff_clk_24_8  VGND ff_rc m=4
xf_24_9  ff_24_9  ff_clk_24_9  VGND ff_rc m=8
xf_24_10 ff_24_10 ff_clk_24_10 VGND ff_rc m=7
xf_25_0  ff_25_0  ff_clk_25_0  VGND ff_rc m=8
xf_25_1  ff_25_1  ff_clk_25_1  VGND ff_rc m=13
xf_25_2  ff_25_2  ff_clk_25_2  VGND ff_rc m=17
xf_25_3  ff_25_3  ff_clk_25_3  VGND ff_rc m=12
xf_25_4  ff_25_4  ff_clk_25_4  VGND ff_rc m=6
xf_25_5  ff_25_5  ff_clk_25_5  VGND ff_rc m=10
xf_25_6  ff_25_6  ff_clk_25_6  VGND ff_rc m=20
xf_25_7  ff_25_7  ff_clk_25_7  VGND ff_rc m=16
xf_25_8  ff_25_8  ff_clk_25_8  VGND ff_rc m=10
xf_25_9  ff_25_9  ff_clk_25_9  VGND ff_rc m=14
xf_25_10 ff_25_10 ff_clk_25_10 VGND ff_rc m=9
xf_25_11 ff_25_11 ff_clk_25_11 VGND ff_rc m=15
xf_26_0  ff_26_0  ff_clk_26_0  VGND ff_rc m=9
xf_26_1  ff_26_1  ff_clk_26_1  VGND ff_rc m=4
xf_26_2  ff_26_2  ff_clk_26_2  VGND ff_rc m=12
xf_26_3  ff_26_3  ff_clk_26_3  VGND ff_rc m=20
xf_26_4  ff_26_4  ff_clk_26_4  VGND ff_rc m=10
xf_26_5  ff_26_5  ff_clk_26_5  VGND ff_rc m=10
xf_26_6  ff_26_6  ff_clk_26_6  VGND ff_rc m=16
xf_26_7  ff_26_7  ff_clk_26_7  VGND ff_rc m=18
xf_26_8  ff_26_8  ff_clk_26_8  VGND ff_rc m=16
xf_26_9  ff_26_9  ff_clk_26_9  VGND ff_rc m=9
xf_27_0  ff_27_0  ff_clk_27_0  VGND ff_rc m=18
xf_27_1  ff_27_1  ff_clk_27_1  VGND ff_rc m=16
xf_27_2  ff_27_2  ff_clk_27_2  VGND ff_rc m=18
xf_27_3  ff_27_3  ff_clk_27_3  VGND ff_rc m=12
xf_27_4  ff_27_4  ff_clk_27_4  VGND ff_rc m=9
xf_27_5  ff_27_5  ff_clk_27_5  VGND ff_rc m=16
xf_27_6  ff_27_6  ff_clk_27_6  VGND ff_rc m=8
xf_27_7  ff_27_7  ff_clk_27_7  VGND ff_rc m=11
xf_27_8  ff_27_8  ff_clk_27_8  VGND ff_rc m=6
xf_28_0  ff_28_0  ff_clk_28_0  VGND ff_rc m=9
xf_28_1  ff_28_1  ff_clk_28_1  VGND ff_rc m=13
xf_28_2  ff_28_2  ff_clk_28_2  VGND ff_rc m=13
xf_28_3  ff_28_3  ff_clk_28_3  VGND ff_rc m=11
xf_28_4  ff_28_4  ff_clk_28_4  VGND ff_rc m=12
xf_28_5  ff_28_5  ff_clk_28_5  VGND ff_rc m=14
xf_28_6  ff_28_6  ff_clk_28_6  VGND ff_rc m=7
xf_28_7  ff_28_7  ff_clk_28_7  VGND ff_rc m=7
xf_28_8  ff_28_8  ff_clk_28_8  VGND ff_rc m=11
xf_28_9  ff_28_9  ff_clk_28_9  VGND ff_rc m=6
xf_28_10 ff_28_10 ff_clk_28_10 VGND ff_rc m=13
xf_28_11 ff_28_11 ff_clk_28_11 VGND ff_rc m=15
xf_28_12 ff_28_12 ff_clk_28_12 VGND ff_rc m=14
xf_29_0  ff_29_0  ff_clk_29_0  VGND ff_rc m=16
xf_29_1  ff_29_1  ff_clk_29_1  VGND ff_rc m=11
xf_29_2  ff_29_2  ff_clk_29_2  VGND ff_rc m=8
xf_29_3  ff_29_3  ff_clk_29_3  VGND ff_rc m=17
xf_29_4  ff_29_4  ff_clk_29_4  VGND ff_rc m=15
xf_29_5  ff_29_5  ff_clk_29_5  VGND ff_rc m=10
xf_29_6  ff_29_6  ff_clk_29_6  VGND ff_rc m=19
xf_29_7  ff_29_7  ff_clk_29_7  VGND ff_rc m=14
xf_29_8  ff_29_8  ff_clk_29_8  VGND ff_rc m=9
xf_29_9  ff_29_9  ff_clk_29_9  VGND ff_rc m=10
xf_29_10 ff_29_10 ff_clk_29_10 VGND ff_rc m=14
xf_29_11 ff_29_11 ff_clk_29_11 VGND ff_rc m=13
xf_29_12 ff_29_12 ff_clk_29_12 VGND ff_rc m=7
xf_30_0  ff_30_0  ff_clk_30_0  VGND ff_rc m=20
xf_30_1  ff_30_1  ff_clk_30_1  VGND ff_rc m=10
xf_30_2  ff_30_2  ff_clk_30_2  VGND ff_rc m=15
xf_30_3  ff_30_3  ff_clk_30_3  VGND ff_rc m=14
xf_30_4  ff_30_4  ff_clk_30_4  VGND ff_rc m=5
xf_30_5  ff_30_5  ff_clk_30_5  VGND ff_rc m=14
xf_30_6  ff_30_6  ff_clk_30_6  VGND ff_rc m=14
xf_30_7  ff_30_7  ff_clk_30_7  VGND ff_rc m=9
xf_31_0  ff_31_0  ff_clk_31_0  VGND ff_rc m=17
xf_31_1  ff_31_1  ff_clk_31_1  VGND ff_rc m=12
xf_31_2  ff_31_2  ff_clk_31_2  VGND ff_rc m=20
xf_31_3  ff_31_3  ff_clk_31_3  VGND ff_rc m=11
xf_31_4  ff_31_4  ff_clk_31_4  VGND ff_rc m=16
xf_31_5  ff_31_5  ff_clk_31_5  VGND ff_rc m=13
xf_31_6  ff_31_6  ff_clk_31_6  VGND ff_rc m=10
xf_31_7  ff_31_7  ff_clk_31_7  VGND ff_rc m=14
xf_31_8  ff_31_8  ff_clk_31_8  VGND ff_rc m=7
xf_31_9  ff_31_9  ff_clk_31_9  VGND ff_rc m=14
xf_31_10 ff_31_10 ff_clk_31_10 VGND ff_rc m=16
xf_31_11 ff_31_11 ff_clk_31_11 VGND ff_rc m=12
xf_31_12 ff_31_12 ff_clk_31_12 VGND ff_rc m=9

C_0_0 co_i_0_0  VGND 0.9F
C_0_1 co_i_0_1  VGND 0.9F
C_0_2 co_i_0_2  VGND 0.9F
C_0_3 co_i_0_3  VGND 0.9F
C_0_4 co_i_0_4  VGND 0.9F
C_0_5 co_i_0_5  VGND 0.9F
C_0_6 co_i_0_6  VGND 0.9F
C_0_7 co_i_0_7  VGND 0.9F
C_0_8 co_i_0_8  VGND 0.9F
C_1_0 co_i_1_0  VGND 0.9F
C_1_1 co_i_1_1  VGND 0.9F
C_1_2 co_i_1_2  VGND 0.9F
C_1_3 co_i_1_3  VGND 0.9F
C_1_4 co_i_1_4  VGND 0.9F
C_1_5 co_i_1_5  VGND 0.9F
C_1_6 co_i_1_6  VGND 0.9F
C_1_7 co_i_1_7  VGND 0.9F
C_1_8 co_i_1_8  VGND 0.9F
C_1_9 co_i_1_9  VGND 0.9F
C_1_10 co_i_1_10 VGND 0.9F
C_2_0 co_i_2_0  VGND 0.9F
C_2_1 co_i_2_1  VGND 0.9F
C_2_2 co_i_2_2  VGND 0.9F
C_2_3 co_i_2_3  VGND 0.9F
C_2_4 co_i_2_4  VGND 0.9F
C_2_5 co_i_2_5  VGND 0.9F
C_2_6 co_i_2_6  VGND 0.9F
C_2_7 co_i_2_7  VGND 0.9F
C_3_0 co_i_3_0  VGND 0.9F
C_3_1 co_i_3_1  VGND 0.9F
C_3_2 co_i_3_2  VGND 0.9F
C_3_3 co_i_3_3  VGND 0.9F
C_3_4 co_i_3_4  VGND 0.9F
C_3_5 co_i_3_5  VGND 0.9F
C_3_6 co_i_3_6  VGND 0.9F
C_3_7 co_i_3_7  VGND 0.9F
C_4_0 co_i_4_0  VGND 0.9F
C_4_1 co_i_4_1  VGND 0.9F
C_4_2 co_i_4_2  VGND 0.9F
C_4_3 co_i_4_3  VGND 0.9F
C_4_4 co_i_4_4  VGND 0.9F
C_4_5 co_i_4_5  VGND 0.9F
C_4_6 co_i_4_6  VGND 0.9F
C_4_7 co_i_4_7  VGND 0.9F
C_5_0 co_i_5_0  VGND 0.9F
C_5_1 co_i_5_1  VGND 0.9F
C_5_2 co_i_5_2  VGND 0.9F
C_5_3 co_i_5_3  VGND 0.9F
C_5_4 co_i_5_4  VGND 0.9F
C_5_5 co_i_5_5  VGND 0.9F
C_5_6 co_i_5_6  VGND 0.9F
C_5_7 co_i_5_7  VGND 0.9F
C_5_8 co_i_5_8  VGND 0.9F
C_5_9 co_i_5_9  VGND 0.9F
C_5_10 co_i_5_10 VGND 0.9F
C_5_11 co_i_5_11 VGND 0.9F
C_6_0 co_i_6_0  VGND 0.9F
C_6_1 co_i_6_1  VGND 0.9F
C_6_2 co_i_6_2  VGND 0.9F
C_6_3 co_i_6_3  VGND 0.9F
C_6_4 co_i_6_4  VGND 0.9F
C_6_5 co_i_6_5  VGND 0.9F
C_6_6 co_i_6_6  VGND 0.9F
C_6_7 co_i_6_7  VGND 0.9F
C_6_8 co_i_6_8  VGND 0.9F
C_6_9 co_i_6_9  VGND 0.9F
C_7_0 co_i_7_0  VGND 0.9F
C_7_1 co_i_7_1  VGND 0.9F
C_7_2 co_i_7_2  VGND 0.9F
C_7_3 co_i_7_3  VGND 0.9F
C_7_4 co_i_7_4  VGND 0.9F
C_7_5 co_i_7_5  VGND 0.9F
C_7_6 co_i_7_6  VGND 0.9F
C_7_7 co_i_7_7  VGND 0.9F
C_7_8 co_i_7_8  VGND 0.9F
C_7_9 co_i_7_9  VGND 0.9F
C_7_10 co_i_7_10 VGND 0.9F
C_7_11 co_i_7_11 VGND 0.9F
C_7_12 co_i_7_12 VGND 0.9F
C_7_13 co_i_7_13 VGND 0.9F
C_7_14 co_i_7_14 VGND 0.9F
C_8_0 co_i_8_0  VGND 0.9F
C_8_1 co_i_8_1  VGND 0.9F
C_8_2 co_i_8_2  VGND 0.9F
C_8_3 co_i_8_3  VGND 0.9F
C_9_0 co_i_9_0  VGND 0.9F
C_9_1 co_i_9_1  VGND 0.9F
C_9_2 co_i_9_2  VGND 0.9F
C_9_3 co_i_9_3  VGND 0.9F
C_9_4 co_i_9_4  VGND 0.9F
C_10_0 co_i_10_0  VGND 0.9F
C_10_1 co_i_10_1  VGND 0.9F
C_10_2 co_i_10_2  VGND 0.9F
C_10_3 co_i_10_3  VGND 0.9F
C_10_4 co_i_10_4  VGND 0.9F
C_10_5 co_i_10_5  VGND 0.9F
C_10_6 co_i_10_6  VGND 0.9F
C_11_0 co_i_11_0  VGND 0.9F
C_11_1 co_i_11_1  VGND 0.9F
C_11_2 co_i_11_2  VGND 0.9F
C_11_3 co_i_11_3  VGND 0.9F
C_11_4 co_i_11_4  VGND 0.9F
C_11_5 co_i_11_5  VGND 0.9F
C_11_6 co_i_11_6  VGND 0.9F
C_11_7 co_i_11_7  VGND 0.9F
C_12_0 co_i_12_0  VGND 0.9F
C_12_1 co_i_12_1  VGND 0.9F
C_12_2 co_i_12_2  VGND 0.9F
C_12_3 co_i_12_3  VGND 0.9F
C_12_4 co_i_12_4  VGND 0.9F
C_13_0 co_i_13_0  VGND 0.9F
C_13_1 co_i_13_1  VGND 0.9F
C_13_2 co_i_13_2  VGND 0.9F
C_13_3 co_i_13_3  VGND 0.9F
C_13_4 co_i_13_4  VGND 0.9F
C_13_5 co_i_13_5  VGND 0.9F
C_13_6 co_i_13_6  VGND 0.9F
C_14_0 co_i_14_0  VGND 0.9F
C_14_1 co_i_14_1  VGND 0.9F
C_14_2 co_i_14_2  VGND 0.9F
C_14_3 co_i_14_3  VGND 0.9F
C_14_4 co_i_14_4  VGND 0.9F
C_15_0 co_i_15_0  VGND 0.9F
C_15_1 co_i_15_1  VGND 0.9F
C_15_2 co_i_15_2  VGND 0.9F
C_15_3 co_i_15_3  VGND 0.9F
C_15_4 co_i_15_4  VGND 0.9F
C_15_5 co_i_15_5  VGND 0.9F
C_15_6 co_i_15_6  VGND 0.9F
C_16_0 co_i_16_0  VGND 0.9F
C_16_1 co_i_16_1  VGND 0.9F
C_16_2 co_i_16_2  VGND 0.9F
C_16_3 co_i_16_3  VGND 0.9F
C_16_4 co_i_16_4  VGND 0.9F
C_16_5 co_i_16_5  VGND 0.9F
C_16_6 co_i_16_6  VGND 0.9F
C_16_7 co_i_16_7  VGND 0.9F
C_16_8 co_i_16_8  VGND 0.9F
C_16_9 co_i_16_9  VGND 0.9F
C_16_10 co_i_16_10 VGND 0.9F
C_17_0 co_i_17_0  VGND 0.9F
C_17_1 co_i_17_1  VGND 0.9F
C_17_2 co_i_17_2  VGND 0.9F
C_17_3 co_i_17_3  VGND 0.9F
C_17_4 co_i_17_4  VGND 0.9F
C_17_5 co_i_17_5  VGND 0.9F
C_17_6 co_i_17_6  VGND 0.9F
C_17_7 co_i_17_7  VGND 0.9F
C_17_8 co_i_17_8  VGND 0.9F
C_17_9 co_i_17_9  VGND 0.9F
C_17_10 co_i_17_10 VGND 0.9F
C_17_11 co_i_17_11 VGND 0.9F
C_17_12 co_i_17_12 VGND 0.9F
C_17_13 co_i_17_13 VGND 0.9F
C_18_0 co_i_18_0  VGND 0.9F
C_18_1 co_i_18_1  VGND 0.9F
C_18_2 co_i_18_2  VGND 0.9F
C_18_3 co_i_18_3  VGND 0.9F
C_18_4 co_i_18_4  VGND 0.9F
C_18_5 co_i_18_5  VGND 0.9F
C_18_6 co_i_18_6  VGND 0.9F
C_18_7 co_i_18_7  VGND 0.9F
C_18_8 co_i_18_8  VGND 0.9F
C_18_9 co_i_18_9  VGND 0.9F
C_18_10 co_i_18_10 VGND 0.9F
C_18_11 co_i_18_11 VGND 0.9F
C_18_12 co_i_18_12 VGND 0.9F
C_19_0 co_i_19_0  VGND 0.9F
C_19_1 co_i_19_1  VGND 0.9F
C_19_2 co_i_19_2  VGND 0.9F
C_19_3 co_i_19_3  VGND 0.9F
C_19_4 co_i_19_4  VGND 0.9F
C_19_5 co_i_19_5  VGND 0.9F
C_19_6 co_i_19_6  VGND 0.9F
C_19_7 co_i_19_7  VGND 0.9F
C_20_0 co_i_20_0  VGND 0.9F
C_20_1 co_i_20_1  VGND 0.9F
C_20_2 co_i_20_2  VGND 0.9F
C_20_3 co_i_20_3  VGND 0.9F
C_20_4 co_i_20_4  VGND 0.9F
C_20_5 co_i_20_5  VGND 0.9F
C_20_6 co_i_20_6  VGND 0.9F
C_20_7 co_i_20_7  VGND 0.9F
C_20_8 co_i_20_8  VGND 0.9F
C_20_9 co_i_20_9  VGND 0.9F
C_20_10 co_i_20_10 VGND 0.9F
C_20_11 co_i_20_11 VGND 0.9F
C_20_12 co_i_20_12 VGND 0.9F
C_20_13 co_i_20_13 VGND 0.9F
C_20_14 co_i_20_14 VGND 0.9F
C_21_0 co_i_21_0  VGND 0.9F
C_21_1 co_i_21_1  VGND 0.9F
C_21_2 co_i_21_2  VGND 0.9F
C_21_3 co_i_21_3  VGND 0.9F
C_21_4 co_i_21_4  VGND 0.9F
C_21_5 co_i_21_5  VGND 0.9F
C_21_6 co_i_21_6  VGND 0.9F
C_21_7 co_i_21_7  VGND 0.9F
C_21_8 co_i_21_8  VGND 0.9F
C_21_9 co_i_21_9  VGND 0.9F
C_21_10 co_i_21_10 VGND 0.9F
C_21_11 co_i_21_11 VGND 0.9F
C_21_12 co_i_21_12 VGND 0.9F
C_22_0 co_i_22_0  VGND 0.9F
C_22_1 co_i_22_1  VGND 0.9F
C_22_2 co_i_22_2  VGND 0.9F
C_22_3 co_i_22_3  VGND 0.9F
C_22_4 co_i_22_4  VGND 0.9F
C_22_5 co_i_22_5  VGND 0.9F
C_22_6 co_i_22_6  VGND 0.9F
C_22_7 co_i_22_7  VGND 0.9F
C_22_8 co_i_22_8  VGND 0.9F
C_22_9 co_i_22_9  VGND 0.9F
C_23_0 co_i_23_0  VGND 0.9F
C_23_1 co_i_23_1  VGND 0.9F
C_23_2 co_i_23_2  VGND 0.9F
C_23_3 co_i_23_3  VGND 0.9F
C_23_4 co_i_23_4  VGND 0.9F
C_23_5 co_i_23_5  VGND 0.9F
C_23_6 co_i_23_6  VGND 0.9F
C_23_7 co_i_23_7  VGND 0.9F
C_23_8 co_i_23_8  VGND 0.9F
C_23_9 co_i_23_9  VGND 0.9F
C_23_10 co_i_23_10 VGND 0.9F
C_23_11 co_i_23_11 VGND 0.9F
C_23_12 co_i_23_12 VGND 0.9F
C_23_13 co_i_23_13 VGND 0.9F
C_23_14 co_i_23_14 VGND 0.9F
C_23_15 co_i_23_15 VGND 0.9F
C_24_0 co_i_24_0  VGND 0.9F
C_24_1 co_i_24_1  VGND 0.9F
C_24_2 co_i_24_2  VGND 0.9F
C_24_3 co_i_24_3  VGND 0.9F
C_24_4 co_i_24_4  VGND 0.9F
C_24_5 co_i_24_5  VGND 0.9F
C_24_6 co_i_24_6  VGND 0.9F
C_24_7 co_i_24_7  VGND 0.9F
C_24_8 co_i_24_8  VGND 0.9F
C_24_9 co_i_24_9  VGND 0.9F
C_24_10 co_i_24_10 VGND 0.9F
C_25_0 co_i_25_0  VGND 0.9F
C_25_1 co_i_25_1  VGND 0.9F
C_25_2 co_i_25_2  VGND 0.9F
C_25_3 co_i_25_3  VGND 0.9F
C_25_4 co_i_25_4  VGND 0.9F
C_25_5 co_i_25_5  VGND 0.9F
C_25_6 co_i_25_6  VGND 0.9F
C_25_7 co_i_25_7  VGND 0.9F
C_25_8 co_i_25_8  VGND 0.9F
C_25_9 co_i_25_9  VGND 0.9F
C_25_10 co_i_25_10 VGND 0.9F
C_25_11 co_i_25_11 VGND 0.9F
C_26_0 co_i_26_0  VGND 0.9F
C_26_1 co_i_26_1  VGND 0.9F
C_26_2 co_i_26_2  VGND 0.9F
C_26_3 co_i_26_3  VGND 0.9F
C_26_4 co_i_26_4  VGND 0.9F
C_26_5 co_i_26_5  VGND 0.9F
C_26_6 co_i_26_6  VGND 0.9F
C_26_7 co_i_26_7  VGND 0.9F
C_26_8 co_i_26_8  VGND 0.9F
C_26_9 co_i_26_9  VGND 0.9F
C_27_0 co_i_27_0  VGND 0.9F
C_27_1 co_i_27_1  VGND 0.9F
C_27_2 co_i_27_2  VGND 0.9F
C_27_3 co_i_27_3  VGND 0.9F
C_27_4 co_i_27_4  VGND 0.9F
C_27_5 co_i_27_5  VGND 0.9F
C_27_6 co_i_27_6  VGND 0.9F
C_27_7 co_i_27_7  VGND 0.9F
C_27_8 co_i_27_8  VGND 0.9F
C_28_0 co_i_28_0  VGND 0.9F
C_28_1 co_i_28_1  VGND 0.9F
C_28_2 co_i_28_2  VGND 0.9F
C_28_3 co_i_28_3  VGND 0.9F
C_28_4 co_i_28_4  VGND 0.9F
C_28_5 co_i_28_5  VGND 0.9F
C_28_6 co_i_28_6  VGND 0.9F
C_28_7 co_i_28_7  VGND 0.9F
C_28_8 co_i_28_8  VGND 0.9F
C_28_9 co_i_28_9  VGND 0.9F
C_28_10 co_i_28_10 VGND 0.9F
C_28_11 co_i_28_11 VGND 0.9F
C_28_12 co_i_28_12 VGND 0.9F
C_29_0 co_i_29_0  VGND 0.9F
C_29_1 co_i_29_1  VGND 0.9F
C_29_2 co_i_29_2  VGND 0.9F
C_29_3 co_i_29_3  VGND 0.9F
C_29_4 co_i_29_4  VGND 0.9F
C_29_5 co_i_29_5  VGND 0.9F
C_29_6 co_i_29_6  VGND 0.9F
C_29_7 co_i_29_7  VGND 0.9F
C_29_8 co_i_29_8  VGND 0.9F
C_29_9 co_i_29_9  VGND 0.9F
C_29_10 co_i_29_10 VGND 0.9F
C_29_11 co_i_29_11 VGND 0.9F
C_29_12 co_i_29_12 VGND 0.9F
C_30_0 co_i_30_0  VGND 0.9F
C_30_1 co_i_30_1  VGND 0.9F
C_30_2 co_i_30_2  VGND 0.9F
C_30_3 co_i_30_3  VGND 0.9F
C_30_4 co_i_30_4  VGND 0.9F
C_30_5 co_i_30_5  VGND 0.9F
C_30_6 co_i_30_6  VGND 0.9F
C_30_7 co_i_30_7  VGND 0.9F
C_31_0 co_i_31_0  VGND 0.9F
C_31_1 co_i_31_1  VGND 0.9F
C_31_2 co_i_31_2  VGND 0.9F
C_31_3 co_i_31_3  VGND 0.9F
C_31_4 co_i_31_4  VGND 0.9F
C_31_5 co_i_31_5  VGND 0.9F
C_31_6 co_i_31_6  VGND 0.9F
C_31_7 co_i_31_7  VGND 0.9F
C_31_8 co_i_31_8  VGND 0.9F
C_31_9 co_i_31_9  VGND 0.9F
C_31_10 co_i_31_10 VGND 0.9F
C_31_11 co_i_31_11 VGND 0.9F
C_31_12 co_i_31_12 VGND 0.9F


.lib     ../../../pdks/sky130A-1.0.227.01/libs.tech/ngspice/sky130.lib.spice ${CORNER}
.include ../../../pdks/sky130A-1.0.227.01/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.include ../../subckts.spice

.temp ${TEMP}
.save all
.tran 0.1n 50n

.end

* NGSPICE file created from sky130_ef_sc_hd__decap_12.ext - technology: sky130A

.subckt sky130_ef_sc_hd__decap_12 VPWR VPB VGND VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
C0 VPWR VGND 2.57fF
.ends


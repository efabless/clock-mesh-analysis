magic
tech sky130A
magscale 1 2
timestamp 1633016303
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 0 -17 672 17
<< locali >>
rect 313 422 408 751
rect 313 388 429 422
rect 25 301 171 367
rect 213 301 359 352
rect 395 325 429 388
rect 465 361 647 424
rect 395 291 564 325
rect 498 99 564 291
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 18 735 208 751
rect 18 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 208 735
rect 18 435 208 701
rect 444 735 634 751
rect 444 701 450 735
rect 484 701 522 735
rect 556 701 594 735
rect 628 701 634 735
rect 444 460 634 701
rect 26 255 92 265
rect 26 221 408 255
rect 26 99 92 221
rect 128 113 306 185
rect 162 79 200 113
rect 234 79 272 113
rect 342 99 408 221
rect 128 73 306 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 24 701 58 735
rect 96 701 130 735
rect 168 701 202 735
rect 450 701 484 735
rect 522 701 556 735
rect 594 701 628 735
rect 128 79 162 113
rect 200 79 234 113
rect 272 79 306 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 450 735
rect 484 701 522 735
rect 556 701 594 735
rect 628 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 128 113
rect 162 79 200 113
rect 234 79 272 113
rect 306 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel locali s 25 301 171 367 6 A1
port 1 nsew signal input
rlabel locali s 213 301 359 352 6 A2
port 2 nsew signal input
rlabel locali s 465 361 647 424 6 B1
port 3 nsew signal input
rlabel locali s 498 99 564 291 6 Y
port 8 nsew signal output
rlabel locali s 395 325 429 388 6 Y
port 8 nsew signal output
rlabel locali s 395 291 564 325 6 Y
port 8 nsew signal output
rlabel locali s 313 422 408 751 6 Y
port 8 nsew signal output
rlabel locali s 313 388 429 422 6 Y
port 8 nsew signal output
rlabel metal1 s 0 51 672 125 6 VGND
port 4 nsew ground bidirectional
rlabel pwell s 0 -17 672 17 8 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 -23 672 23 8 VNB
port 5 nsew ground bidirectional
rlabel nwell s -66 377 738 897 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 791 672 837 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 689 672 763 6 VPWR
port 7 nsew power bidirectional
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 672 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 286066
string GDS_START 277112
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1633016076
<< checkpaint >>
rect -1260 -1260 2142 2648
<< nwell >>
rect 0 0 882 1388
<< pmos >>
rect 171 189 201 1199
rect 257 189 307 1199
rect 363 189 413 1199
rect 469 189 519 1199
rect 575 189 625 1199
rect 681 189 711 1199
<< pdiff >>
rect 111 1187 171 1199
rect 111 1153 126 1187
rect 160 1153 171 1187
rect 111 1119 171 1153
rect 111 1085 126 1119
rect 160 1085 171 1119
rect 111 1051 171 1085
rect 111 1017 126 1051
rect 160 1017 171 1051
rect 111 983 171 1017
rect 111 949 126 983
rect 160 949 171 983
rect 111 915 171 949
rect 111 881 126 915
rect 160 881 171 915
rect 111 847 171 881
rect 111 813 126 847
rect 160 813 171 847
rect 111 779 171 813
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 1187 257 1199
rect 201 1153 212 1187
rect 246 1153 257 1187
rect 201 1119 257 1153
rect 201 1085 212 1119
rect 246 1085 257 1119
rect 201 1051 257 1085
rect 201 1017 212 1051
rect 246 1017 257 1051
rect 201 983 257 1017
rect 201 949 212 983
rect 246 949 257 983
rect 201 915 257 949
rect 201 881 212 915
rect 246 881 257 915
rect 201 847 257 881
rect 201 813 212 847
rect 246 813 257 847
rect 201 779 257 813
rect 201 745 212 779
rect 246 745 257 779
rect 201 711 257 745
rect 201 677 212 711
rect 246 677 257 711
rect 201 643 257 677
rect 201 609 212 643
rect 246 609 257 643
rect 201 575 257 609
rect 201 541 212 575
rect 246 541 257 575
rect 201 507 257 541
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 307 1187 363 1199
rect 307 1153 318 1187
rect 352 1153 363 1187
rect 307 1119 363 1153
rect 307 1085 318 1119
rect 352 1085 363 1119
rect 307 1051 363 1085
rect 307 1017 318 1051
rect 352 1017 363 1051
rect 307 983 363 1017
rect 307 949 318 983
rect 352 949 363 983
rect 307 915 363 949
rect 307 881 318 915
rect 352 881 363 915
rect 307 847 363 881
rect 307 813 318 847
rect 352 813 363 847
rect 307 779 363 813
rect 307 745 318 779
rect 352 745 363 779
rect 307 711 363 745
rect 307 677 318 711
rect 352 677 363 711
rect 307 643 363 677
rect 307 609 318 643
rect 352 609 363 643
rect 307 575 363 609
rect 307 541 318 575
rect 352 541 363 575
rect 307 507 363 541
rect 307 473 318 507
rect 352 473 363 507
rect 307 439 363 473
rect 307 405 318 439
rect 352 405 363 439
rect 307 371 363 405
rect 307 337 318 371
rect 352 337 363 371
rect 307 303 363 337
rect 307 269 318 303
rect 352 269 363 303
rect 307 235 363 269
rect 307 201 318 235
rect 352 201 363 235
rect 307 189 363 201
rect 413 1187 469 1199
rect 413 1153 424 1187
rect 458 1153 469 1187
rect 413 1119 469 1153
rect 413 1085 424 1119
rect 458 1085 469 1119
rect 413 1051 469 1085
rect 413 1017 424 1051
rect 458 1017 469 1051
rect 413 983 469 1017
rect 413 949 424 983
rect 458 949 469 983
rect 413 915 469 949
rect 413 881 424 915
rect 458 881 469 915
rect 413 847 469 881
rect 413 813 424 847
rect 458 813 469 847
rect 413 779 469 813
rect 413 745 424 779
rect 458 745 469 779
rect 413 711 469 745
rect 413 677 424 711
rect 458 677 469 711
rect 413 643 469 677
rect 413 609 424 643
rect 458 609 469 643
rect 413 575 469 609
rect 413 541 424 575
rect 458 541 469 575
rect 413 507 469 541
rect 413 473 424 507
rect 458 473 469 507
rect 413 439 469 473
rect 413 405 424 439
rect 458 405 469 439
rect 413 371 469 405
rect 413 337 424 371
rect 458 337 469 371
rect 413 303 469 337
rect 413 269 424 303
rect 458 269 469 303
rect 413 235 469 269
rect 413 201 424 235
rect 458 201 469 235
rect 413 189 469 201
rect 519 1187 575 1199
rect 519 1153 530 1187
rect 564 1153 575 1187
rect 519 1119 575 1153
rect 519 1085 530 1119
rect 564 1085 575 1119
rect 519 1051 575 1085
rect 519 1017 530 1051
rect 564 1017 575 1051
rect 519 983 575 1017
rect 519 949 530 983
rect 564 949 575 983
rect 519 915 575 949
rect 519 881 530 915
rect 564 881 575 915
rect 519 847 575 881
rect 519 813 530 847
rect 564 813 575 847
rect 519 779 575 813
rect 519 745 530 779
rect 564 745 575 779
rect 519 711 575 745
rect 519 677 530 711
rect 564 677 575 711
rect 519 643 575 677
rect 519 609 530 643
rect 564 609 575 643
rect 519 575 575 609
rect 519 541 530 575
rect 564 541 575 575
rect 519 507 575 541
rect 519 473 530 507
rect 564 473 575 507
rect 519 439 575 473
rect 519 405 530 439
rect 564 405 575 439
rect 519 371 575 405
rect 519 337 530 371
rect 564 337 575 371
rect 519 303 575 337
rect 519 269 530 303
rect 564 269 575 303
rect 519 235 575 269
rect 519 201 530 235
rect 564 201 575 235
rect 519 189 575 201
rect 625 1187 681 1199
rect 625 1153 636 1187
rect 670 1153 681 1187
rect 625 1119 681 1153
rect 625 1085 636 1119
rect 670 1085 681 1119
rect 625 1051 681 1085
rect 625 1017 636 1051
rect 670 1017 681 1051
rect 625 983 681 1017
rect 625 949 636 983
rect 670 949 681 983
rect 625 915 681 949
rect 625 881 636 915
rect 670 881 681 915
rect 625 847 681 881
rect 625 813 636 847
rect 670 813 681 847
rect 625 779 681 813
rect 625 745 636 779
rect 670 745 681 779
rect 625 711 681 745
rect 625 677 636 711
rect 670 677 681 711
rect 625 643 681 677
rect 625 609 636 643
rect 670 609 681 643
rect 625 575 681 609
rect 625 541 636 575
rect 670 541 681 575
rect 625 507 681 541
rect 625 473 636 507
rect 670 473 681 507
rect 625 439 681 473
rect 625 405 636 439
rect 670 405 681 439
rect 625 371 681 405
rect 625 337 636 371
rect 670 337 681 371
rect 625 303 681 337
rect 625 269 636 303
rect 670 269 681 303
rect 625 235 681 269
rect 625 201 636 235
rect 670 201 681 235
rect 625 189 681 201
rect 711 1187 771 1199
rect 711 1153 722 1187
rect 756 1153 771 1187
rect 711 1119 771 1153
rect 711 1085 722 1119
rect 756 1085 771 1119
rect 711 1051 771 1085
rect 711 1017 722 1051
rect 756 1017 771 1051
rect 711 983 771 1017
rect 711 949 722 983
rect 756 949 771 983
rect 711 915 771 949
rect 711 881 722 915
rect 756 881 771 915
rect 711 847 771 881
rect 711 813 722 847
rect 756 813 771 847
rect 711 779 771 813
rect 711 745 722 779
rect 756 745 771 779
rect 711 711 771 745
rect 711 677 722 711
rect 756 677 771 711
rect 711 643 771 677
rect 711 609 722 643
rect 756 609 771 643
rect 711 575 771 609
rect 711 541 722 575
rect 756 541 771 575
rect 711 507 771 541
rect 711 473 722 507
rect 756 473 771 507
rect 711 439 771 473
rect 711 405 722 439
rect 756 405 771 439
rect 711 371 771 405
rect 711 337 722 371
rect 756 337 771 371
rect 711 303 771 337
rect 711 269 722 303
rect 756 269 771 303
rect 711 235 771 269
rect 711 201 722 235
rect 756 201 771 235
rect 711 189 771 201
<< pdiffc >>
rect 126 1153 160 1187
rect 126 1085 160 1119
rect 126 1017 160 1051
rect 126 949 160 983
rect 126 881 160 915
rect 126 813 160 847
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 1153 246 1187
rect 212 1085 246 1119
rect 212 1017 246 1051
rect 212 949 246 983
rect 212 881 246 915
rect 212 813 246 847
rect 212 745 246 779
rect 212 677 246 711
rect 212 609 246 643
rect 212 541 246 575
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 318 1153 352 1187
rect 318 1085 352 1119
rect 318 1017 352 1051
rect 318 949 352 983
rect 318 881 352 915
rect 318 813 352 847
rect 318 745 352 779
rect 318 677 352 711
rect 318 609 352 643
rect 318 541 352 575
rect 318 473 352 507
rect 318 405 352 439
rect 318 337 352 371
rect 318 269 352 303
rect 318 201 352 235
rect 424 1153 458 1187
rect 424 1085 458 1119
rect 424 1017 458 1051
rect 424 949 458 983
rect 424 881 458 915
rect 424 813 458 847
rect 424 745 458 779
rect 424 677 458 711
rect 424 609 458 643
rect 424 541 458 575
rect 424 473 458 507
rect 424 405 458 439
rect 424 337 458 371
rect 424 269 458 303
rect 424 201 458 235
rect 530 1153 564 1187
rect 530 1085 564 1119
rect 530 1017 564 1051
rect 530 949 564 983
rect 530 881 564 915
rect 530 813 564 847
rect 530 745 564 779
rect 530 677 564 711
rect 530 609 564 643
rect 530 541 564 575
rect 530 473 564 507
rect 530 405 564 439
rect 530 337 564 371
rect 530 269 564 303
rect 530 201 564 235
rect 636 1153 670 1187
rect 636 1085 670 1119
rect 636 1017 670 1051
rect 636 949 670 983
rect 636 881 670 915
rect 636 813 670 847
rect 636 745 670 779
rect 636 677 670 711
rect 636 609 670 643
rect 636 541 670 575
rect 636 473 670 507
rect 636 405 670 439
rect 636 337 670 371
rect 636 269 670 303
rect 636 201 670 235
rect 722 1153 756 1187
rect 722 1085 756 1119
rect 722 1017 756 1051
rect 722 949 756 983
rect 722 881 756 915
rect 722 813 756 847
rect 722 745 756 779
rect 722 677 756 711
rect 722 609 756 643
rect 722 541 756 575
rect 722 473 756 507
rect 722 405 756 439
rect 722 337 756 371
rect 722 269 756 303
rect 722 201 756 235
<< nsubdiff >>
rect 41 1187 111 1199
rect 41 1153 58 1187
rect 92 1153 111 1187
rect 41 1119 111 1153
rect 41 1085 58 1119
rect 92 1085 111 1119
rect 41 1051 111 1085
rect 41 1017 58 1051
rect 92 1017 111 1051
rect 41 983 111 1017
rect 41 949 58 983
rect 92 949 111 983
rect 41 915 111 949
rect 41 881 58 915
rect 92 881 111 915
rect 41 847 111 881
rect 41 813 58 847
rect 92 813 111 847
rect 41 779 111 813
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 771 1187 841 1199
rect 771 1153 790 1187
rect 824 1153 841 1187
rect 771 1119 841 1153
rect 771 1085 790 1119
rect 824 1085 841 1119
rect 771 1051 841 1085
rect 771 1017 790 1051
rect 824 1017 841 1051
rect 771 983 841 1017
rect 771 949 790 983
rect 824 949 841 983
rect 771 915 841 949
rect 771 881 790 915
rect 824 881 841 915
rect 771 847 841 881
rect 771 813 790 847
rect 824 813 841 847
rect 771 779 841 813
rect 771 745 790 779
rect 824 745 841 779
rect 771 711 841 745
rect 771 677 790 711
rect 824 677 841 711
rect 771 643 841 677
rect 771 609 790 643
rect 824 609 841 643
rect 771 575 841 609
rect 771 541 790 575
rect 824 541 841 575
rect 771 507 841 541
rect 771 473 790 507
rect 824 473 841 507
rect 771 439 841 473
rect 771 405 790 439
rect 824 405 841 439
rect 771 371 841 405
rect 771 337 790 371
rect 824 337 841 371
rect 771 303 841 337
rect 771 269 790 303
rect 824 269 841 303
rect 771 235 841 269
rect 771 201 790 235
rect 824 201 841 235
rect 771 189 841 201
<< nsubdiffcont >>
rect 58 1153 92 1187
rect 58 1085 92 1119
rect 58 1017 92 1051
rect 58 949 92 983
rect 58 881 92 915
rect 58 813 92 847
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 790 1153 824 1187
rect 790 1085 824 1119
rect 790 1017 824 1051
rect 790 949 824 983
rect 790 881 824 915
rect 790 813 824 847
rect 790 745 824 779
rect 790 677 824 711
rect 790 609 824 643
rect 790 541 824 575
rect 790 473 824 507
rect 790 405 824 439
rect 790 337 824 371
rect 790 269 824 303
rect 790 201 824 235
<< poly >>
rect 243 1367 639 1388
rect 120 1281 201 1297
rect 120 1247 136 1281
rect 170 1247 201 1281
rect 243 1265 288 1367
rect 594 1265 639 1367
rect 243 1249 639 1265
rect 681 1281 762 1297
rect 120 1231 201 1247
rect 171 1199 201 1231
rect 257 1199 307 1249
rect 363 1199 413 1249
rect 469 1199 519 1249
rect 575 1199 625 1249
rect 681 1247 712 1281
rect 746 1247 762 1281
rect 681 1231 762 1247
rect 681 1199 711 1231
rect 171 157 201 189
rect 120 141 201 157
rect 120 107 136 141
rect 170 107 201 141
rect 257 139 307 189
rect 363 139 413 189
rect 469 139 519 189
rect 575 139 625 189
rect 681 157 711 189
rect 681 141 762 157
rect 120 91 201 107
rect 243 123 639 139
rect 243 21 288 123
rect 594 21 639 123
rect 681 107 712 141
rect 746 107 762 141
rect 681 91 762 107
rect 243 0 639 21
<< polycont >>
rect 136 1247 170 1281
rect 288 1265 594 1367
rect 712 1247 746 1281
rect 136 107 170 141
rect 288 21 594 123
rect 712 107 746 141
<< locali >>
rect 266 1369 616 1388
rect 120 1281 186 1297
rect 120 1247 136 1281
rect 170 1247 186 1281
rect 266 1263 280 1369
rect 602 1263 616 1369
rect 266 1249 616 1263
rect 696 1281 762 1297
rect 120 1231 186 1247
rect 696 1247 712 1281
rect 746 1247 762 1281
rect 696 1231 762 1247
rect 120 1203 160 1231
rect 722 1203 762 1231
rect 41 1187 160 1203
rect 41 1153 58 1187
rect 92 1179 126 1187
rect 94 1153 126 1179
rect 41 1145 60 1153
rect 94 1145 160 1153
rect 41 1119 160 1145
rect 41 1085 58 1119
rect 92 1107 126 1119
rect 94 1085 126 1107
rect 41 1073 60 1085
rect 94 1073 160 1085
rect 41 1051 160 1073
rect 41 1017 58 1051
rect 92 1035 126 1051
rect 94 1017 126 1035
rect 41 1001 60 1017
rect 94 1001 160 1017
rect 41 983 160 1001
rect 41 949 58 983
rect 92 963 126 983
rect 94 949 126 963
rect 41 929 60 949
rect 94 929 160 949
rect 41 915 160 929
rect 41 881 58 915
rect 92 891 126 915
rect 94 881 126 891
rect 41 857 60 881
rect 94 857 160 881
rect 41 847 160 857
rect 41 813 58 847
rect 92 819 126 847
rect 94 813 126 819
rect 41 785 60 813
rect 94 785 160 813
rect 41 779 160 785
rect 41 745 58 779
rect 92 747 126 779
rect 94 745 126 747
rect 41 713 60 745
rect 94 713 160 745
rect 41 711 160 713
rect 41 677 58 711
rect 92 677 126 711
rect 41 675 160 677
rect 41 643 60 675
rect 94 643 160 675
rect 41 609 58 643
rect 94 641 126 643
rect 92 609 126 641
rect 41 603 160 609
rect 41 575 60 603
rect 94 575 160 603
rect 41 541 58 575
rect 94 569 126 575
rect 92 541 126 569
rect 41 531 160 541
rect 41 507 60 531
rect 94 507 160 531
rect 41 473 58 507
rect 94 497 126 507
rect 92 473 126 497
rect 41 459 160 473
rect 41 439 60 459
rect 94 439 160 459
rect 41 405 58 439
rect 94 425 126 439
rect 92 405 126 425
rect 41 387 160 405
rect 41 371 60 387
rect 94 371 160 387
rect 41 337 58 371
rect 94 353 126 371
rect 92 337 126 353
rect 41 315 160 337
rect 41 303 60 315
rect 94 303 160 315
rect 41 269 58 303
rect 94 281 126 303
rect 92 269 126 281
rect 41 243 160 269
rect 41 235 60 243
rect 94 235 160 243
rect 41 201 58 235
rect 94 209 126 235
rect 92 201 126 209
rect 41 185 160 201
rect 212 1187 246 1203
rect 212 1119 246 1145
rect 212 1051 246 1073
rect 212 983 246 1001
rect 212 915 246 929
rect 212 847 246 857
rect 212 779 246 785
rect 212 711 246 713
rect 212 675 246 677
rect 212 603 246 609
rect 212 531 246 541
rect 212 459 246 473
rect 212 387 246 405
rect 212 315 246 337
rect 212 243 246 269
rect 212 185 246 201
rect 318 1187 352 1203
rect 318 1119 352 1145
rect 318 1051 352 1073
rect 318 983 352 1001
rect 318 915 352 929
rect 318 847 352 857
rect 318 779 352 785
rect 318 711 352 713
rect 318 675 352 677
rect 318 603 352 609
rect 318 531 352 541
rect 318 459 352 473
rect 318 387 352 405
rect 318 315 352 337
rect 318 243 352 269
rect 318 185 352 201
rect 424 1187 458 1203
rect 424 1119 458 1145
rect 424 1051 458 1073
rect 424 983 458 1001
rect 424 915 458 929
rect 424 847 458 857
rect 424 779 458 785
rect 424 711 458 713
rect 424 675 458 677
rect 424 603 458 609
rect 424 531 458 541
rect 424 459 458 473
rect 424 387 458 405
rect 424 315 458 337
rect 424 243 458 269
rect 424 185 458 201
rect 530 1187 564 1203
rect 530 1119 564 1145
rect 530 1051 564 1073
rect 530 983 564 1001
rect 530 915 564 929
rect 530 847 564 857
rect 530 779 564 785
rect 530 711 564 713
rect 530 675 564 677
rect 530 603 564 609
rect 530 531 564 541
rect 530 459 564 473
rect 530 387 564 405
rect 530 315 564 337
rect 530 243 564 269
rect 530 185 564 201
rect 636 1187 670 1203
rect 636 1119 670 1145
rect 636 1051 670 1073
rect 636 983 670 1001
rect 636 915 670 929
rect 636 847 670 857
rect 636 779 670 785
rect 636 711 670 713
rect 636 675 670 677
rect 636 603 670 609
rect 636 531 670 541
rect 636 459 670 473
rect 636 387 670 405
rect 636 315 670 337
rect 636 243 670 269
rect 636 185 670 201
rect 722 1187 841 1203
rect 756 1179 790 1187
rect 756 1153 788 1179
rect 824 1153 841 1187
rect 722 1145 788 1153
rect 822 1145 841 1153
rect 722 1119 841 1145
rect 756 1107 790 1119
rect 756 1085 788 1107
rect 824 1085 841 1119
rect 722 1073 788 1085
rect 822 1073 841 1085
rect 722 1051 841 1073
rect 756 1035 790 1051
rect 756 1017 788 1035
rect 824 1017 841 1051
rect 722 1001 788 1017
rect 822 1001 841 1017
rect 722 983 841 1001
rect 756 963 790 983
rect 756 949 788 963
rect 824 949 841 983
rect 722 929 788 949
rect 822 929 841 949
rect 722 915 841 929
rect 756 891 790 915
rect 756 881 788 891
rect 824 881 841 915
rect 722 857 788 881
rect 822 857 841 881
rect 722 847 841 857
rect 756 819 790 847
rect 756 813 788 819
rect 824 813 841 847
rect 722 785 788 813
rect 822 785 841 813
rect 722 779 841 785
rect 756 747 790 779
rect 756 745 788 747
rect 824 745 841 779
rect 722 713 788 745
rect 822 713 841 745
rect 722 711 841 713
rect 756 677 790 711
rect 824 677 841 711
rect 722 675 841 677
rect 722 643 788 675
rect 822 643 841 675
rect 756 641 788 643
rect 756 609 790 641
rect 824 609 841 643
rect 722 603 841 609
rect 722 575 788 603
rect 822 575 841 603
rect 756 569 788 575
rect 756 541 790 569
rect 824 541 841 575
rect 722 531 841 541
rect 722 507 788 531
rect 822 507 841 531
rect 756 497 788 507
rect 756 473 790 497
rect 824 473 841 507
rect 722 459 841 473
rect 722 439 788 459
rect 822 439 841 459
rect 756 425 788 439
rect 756 405 790 425
rect 824 405 841 439
rect 722 387 841 405
rect 722 371 788 387
rect 822 371 841 387
rect 756 353 788 371
rect 756 337 790 353
rect 824 337 841 371
rect 722 315 841 337
rect 722 303 788 315
rect 822 303 841 315
rect 756 281 788 303
rect 756 269 790 281
rect 824 269 841 303
rect 722 243 841 269
rect 722 235 788 243
rect 822 235 841 243
rect 756 209 788 235
rect 756 201 790 209
rect 824 201 841 235
rect 722 185 841 201
rect 120 157 160 185
rect 722 157 762 185
rect 120 141 186 157
rect 120 107 136 141
rect 170 107 186 141
rect 696 141 762 157
rect 120 91 186 107
rect 266 125 616 139
rect 266 19 280 125
rect 602 19 616 125
rect 696 107 712 141
rect 746 107 762 141
rect 696 91 762 107
rect 266 0 616 19
<< viali >>
rect 280 1367 602 1369
rect 280 1265 288 1367
rect 288 1265 594 1367
rect 594 1265 602 1367
rect 280 1263 602 1265
rect 60 1153 92 1179
rect 92 1153 94 1179
rect 60 1145 94 1153
rect 60 1085 92 1107
rect 92 1085 94 1107
rect 60 1073 94 1085
rect 60 1017 92 1035
rect 92 1017 94 1035
rect 60 1001 94 1017
rect 60 949 92 963
rect 92 949 94 963
rect 60 929 94 949
rect 60 881 92 891
rect 92 881 94 891
rect 60 857 94 881
rect 60 813 92 819
rect 92 813 94 819
rect 60 785 94 813
rect 60 745 92 747
rect 92 745 94 747
rect 60 713 94 745
rect 60 643 94 675
rect 60 641 92 643
rect 92 641 94 643
rect 60 575 94 603
rect 60 569 92 575
rect 92 569 94 575
rect 60 507 94 531
rect 60 497 92 507
rect 92 497 94 507
rect 60 439 94 459
rect 60 425 92 439
rect 92 425 94 439
rect 60 371 94 387
rect 60 353 92 371
rect 92 353 94 371
rect 60 303 94 315
rect 60 281 92 303
rect 92 281 94 303
rect 60 235 94 243
rect 60 209 92 235
rect 92 209 94 235
rect 212 1153 246 1179
rect 212 1145 246 1153
rect 212 1085 246 1107
rect 212 1073 246 1085
rect 212 1017 246 1035
rect 212 1001 246 1017
rect 212 949 246 963
rect 212 929 246 949
rect 212 881 246 891
rect 212 857 246 881
rect 212 813 246 819
rect 212 785 246 813
rect 212 745 246 747
rect 212 713 246 745
rect 212 643 246 675
rect 212 641 246 643
rect 212 575 246 603
rect 212 569 246 575
rect 212 507 246 531
rect 212 497 246 507
rect 212 439 246 459
rect 212 425 246 439
rect 212 371 246 387
rect 212 353 246 371
rect 212 303 246 315
rect 212 281 246 303
rect 212 235 246 243
rect 212 209 246 235
rect 318 1153 352 1179
rect 318 1145 352 1153
rect 318 1085 352 1107
rect 318 1073 352 1085
rect 318 1017 352 1035
rect 318 1001 352 1017
rect 318 949 352 963
rect 318 929 352 949
rect 318 881 352 891
rect 318 857 352 881
rect 318 813 352 819
rect 318 785 352 813
rect 318 745 352 747
rect 318 713 352 745
rect 318 643 352 675
rect 318 641 352 643
rect 318 575 352 603
rect 318 569 352 575
rect 318 507 352 531
rect 318 497 352 507
rect 318 439 352 459
rect 318 425 352 439
rect 318 371 352 387
rect 318 353 352 371
rect 318 303 352 315
rect 318 281 352 303
rect 318 235 352 243
rect 318 209 352 235
rect 424 1153 458 1179
rect 424 1145 458 1153
rect 424 1085 458 1107
rect 424 1073 458 1085
rect 424 1017 458 1035
rect 424 1001 458 1017
rect 424 949 458 963
rect 424 929 458 949
rect 424 881 458 891
rect 424 857 458 881
rect 424 813 458 819
rect 424 785 458 813
rect 424 745 458 747
rect 424 713 458 745
rect 424 643 458 675
rect 424 641 458 643
rect 424 575 458 603
rect 424 569 458 575
rect 424 507 458 531
rect 424 497 458 507
rect 424 439 458 459
rect 424 425 458 439
rect 424 371 458 387
rect 424 353 458 371
rect 424 303 458 315
rect 424 281 458 303
rect 424 235 458 243
rect 424 209 458 235
rect 530 1153 564 1179
rect 530 1145 564 1153
rect 530 1085 564 1107
rect 530 1073 564 1085
rect 530 1017 564 1035
rect 530 1001 564 1017
rect 530 949 564 963
rect 530 929 564 949
rect 530 881 564 891
rect 530 857 564 881
rect 530 813 564 819
rect 530 785 564 813
rect 530 745 564 747
rect 530 713 564 745
rect 530 643 564 675
rect 530 641 564 643
rect 530 575 564 603
rect 530 569 564 575
rect 530 507 564 531
rect 530 497 564 507
rect 530 439 564 459
rect 530 425 564 439
rect 530 371 564 387
rect 530 353 564 371
rect 530 303 564 315
rect 530 281 564 303
rect 530 235 564 243
rect 530 209 564 235
rect 636 1153 670 1179
rect 636 1145 670 1153
rect 636 1085 670 1107
rect 636 1073 670 1085
rect 636 1017 670 1035
rect 636 1001 670 1017
rect 636 949 670 963
rect 636 929 670 949
rect 636 881 670 891
rect 636 857 670 881
rect 636 813 670 819
rect 636 785 670 813
rect 636 745 670 747
rect 636 713 670 745
rect 636 643 670 675
rect 636 641 670 643
rect 636 575 670 603
rect 636 569 670 575
rect 636 507 670 531
rect 636 497 670 507
rect 636 439 670 459
rect 636 425 670 439
rect 636 371 670 387
rect 636 353 670 371
rect 636 303 670 315
rect 636 281 670 303
rect 636 235 670 243
rect 636 209 670 235
rect 788 1153 790 1179
rect 790 1153 822 1179
rect 788 1145 822 1153
rect 788 1085 790 1107
rect 790 1085 822 1107
rect 788 1073 822 1085
rect 788 1017 790 1035
rect 790 1017 822 1035
rect 788 1001 822 1017
rect 788 949 790 963
rect 790 949 822 963
rect 788 929 822 949
rect 788 881 790 891
rect 790 881 822 891
rect 788 857 822 881
rect 788 813 790 819
rect 790 813 822 819
rect 788 785 822 813
rect 788 745 790 747
rect 790 745 822 747
rect 788 713 822 745
rect 788 643 822 675
rect 788 641 790 643
rect 790 641 822 643
rect 788 575 822 603
rect 788 569 790 575
rect 790 569 822 575
rect 788 507 822 531
rect 788 497 790 507
rect 790 497 822 507
rect 788 439 822 459
rect 788 425 790 439
rect 790 425 822 439
rect 788 371 822 387
rect 788 353 790 371
rect 790 353 822 371
rect 788 303 822 315
rect 788 281 790 303
rect 790 281 822 303
rect 788 235 822 243
rect 788 209 790 235
rect 790 209 822 235
rect 280 123 602 125
rect 280 21 288 123
rect 288 21 594 123
rect 594 21 602 123
rect 280 19 602 21
<< metal1 >>
rect 264 1369 618 1388
rect 264 1263 280 1369
rect 602 1263 618 1369
rect 264 1251 618 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 203 1179 255 1191
rect 203 1145 212 1179
rect 246 1145 255 1179
rect 203 1107 255 1145
rect 203 1073 212 1107
rect 246 1073 255 1107
rect 203 1035 255 1073
rect 203 1001 212 1035
rect 246 1001 255 1035
rect 203 963 255 1001
rect 203 929 212 963
rect 246 929 255 963
rect 203 891 255 929
rect 203 857 212 891
rect 246 857 255 891
rect 203 819 255 857
rect 203 785 212 819
rect 246 785 255 819
rect 203 747 255 785
rect 203 713 212 747
rect 246 713 255 747
rect 203 675 255 713
rect 203 641 212 675
rect 246 641 255 675
rect 203 639 255 641
rect 203 575 212 587
rect 246 575 255 587
rect 203 511 212 523
rect 246 511 255 523
rect 203 447 212 459
rect 246 447 255 459
rect 203 387 255 395
rect 203 383 212 387
rect 246 383 255 387
rect 203 319 255 331
rect 203 255 255 267
rect 203 197 255 203
rect 309 1185 361 1191
rect 309 1121 361 1133
rect 309 1057 361 1069
rect 309 1001 318 1005
rect 352 1001 361 1005
rect 309 993 361 1001
rect 309 929 318 941
rect 352 929 361 941
rect 309 865 318 877
rect 352 865 361 877
rect 309 801 318 813
rect 352 801 361 813
rect 309 747 361 749
rect 309 713 318 747
rect 352 713 361 747
rect 309 675 361 713
rect 309 641 318 675
rect 352 641 361 675
rect 309 603 361 641
rect 309 569 318 603
rect 352 569 361 603
rect 309 531 361 569
rect 309 497 318 531
rect 352 497 361 531
rect 309 459 361 497
rect 309 425 318 459
rect 352 425 361 459
rect 309 387 361 425
rect 309 353 318 387
rect 352 353 361 387
rect 309 315 361 353
rect 309 281 318 315
rect 352 281 361 315
rect 309 243 361 281
rect 309 209 318 243
rect 352 209 361 243
rect 309 197 361 209
rect 415 1179 467 1191
rect 415 1145 424 1179
rect 458 1145 467 1179
rect 415 1107 467 1145
rect 415 1073 424 1107
rect 458 1073 467 1107
rect 415 1035 467 1073
rect 415 1001 424 1035
rect 458 1001 467 1035
rect 415 963 467 1001
rect 415 929 424 963
rect 458 929 467 963
rect 415 891 467 929
rect 415 857 424 891
rect 458 857 467 891
rect 415 819 467 857
rect 415 785 424 819
rect 458 785 467 819
rect 415 747 467 785
rect 415 713 424 747
rect 458 713 467 747
rect 415 675 467 713
rect 415 641 424 675
rect 458 641 467 675
rect 415 639 467 641
rect 415 575 424 587
rect 458 575 467 587
rect 415 511 424 523
rect 458 511 467 523
rect 415 447 424 459
rect 458 447 467 459
rect 415 387 467 395
rect 415 383 424 387
rect 458 383 467 387
rect 415 319 467 331
rect 415 255 467 267
rect 415 197 467 203
rect 521 1185 573 1191
rect 521 1121 573 1133
rect 521 1057 573 1069
rect 521 1001 530 1005
rect 564 1001 573 1005
rect 521 993 573 1001
rect 521 929 530 941
rect 564 929 573 941
rect 521 865 530 877
rect 564 865 573 877
rect 521 801 530 813
rect 564 801 573 813
rect 521 747 573 749
rect 521 713 530 747
rect 564 713 573 747
rect 521 675 573 713
rect 521 641 530 675
rect 564 641 573 675
rect 521 603 573 641
rect 521 569 530 603
rect 564 569 573 603
rect 521 531 573 569
rect 521 497 530 531
rect 564 497 573 531
rect 521 459 573 497
rect 521 425 530 459
rect 564 425 573 459
rect 521 387 573 425
rect 521 353 530 387
rect 564 353 573 387
rect 521 315 573 353
rect 521 281 530 315
rect 564 281 573 315
rect 521 243 573 281
rect 521 209 530 243
rect 564 209 573 243
rect 521 197 573 209
rect 627 1179 679 1191
rect 627 1145 636 1179
rect 670 1145 679 1179
rect 627 1107 679 1145
rect 627 1073 636 1107
rect 670 1073 679 1107
rect 627 1035 679 1073
rect 627 1001 636 1035
rect 670 1001 679 1035
rect 627 963 679 1001
rect 627 929 636 963
rect 670 929 679 963
rect 627 891 679 929
rect 627 857 636 891
rect 670 857 679 891
rect 627 819 679 857
rect 627 785 636 819
rect 670 785 679 819
rect 627 747 679 785
rect 627 713 636 747
rect 670 713 679 747
rect 627 675 679 713
rect 627 641 636 675
rect 670 641 679 675
rect 627 639 679 641
rect 627 575 636 587
rect 670 575 679 587
rect 627 511 636 523
rect 670 511 679 523
rect 627 447 636 459
rect 670 447 679 459
rect 627 387 679 395
rect 627 383 636 387
rect 670 383 679 387
rect 627 319 679 331
rect 627 255 679 267
rect 627 197 679 203
rect 782 1179 841 1191
rect 782 1145 788 1179
rect 822 1145 841 1179
rect 782 1107 841 1145
rect 782 1073 788 1107
rect 822 1073 841 1107
rect 782 1035 841 1073
rect 782 1001 788 1035
rect 822 1001 841 1035
rect 782 963 841 1001
rect 782 929 788 963
rect 822 929 841 963
rect 782 891 841 929
rect 782 857 788 891
rect 822 857 841 891
rect 782 819 841 857
rect 782 785 788 819
rect 822 785 841 819
rect 782 747 841 785
rect 782 713 788 747
rect 822 713 841 747
rect 782 675 841 713
rect 782 641 788 675
rect 822 641 841 675
rect 782 603 841 641
rect 782 569 788 603
rect 822 569 841 603
rect 782 531 841 569
rect 782 497 788 531
rect 822 497 841 531
rect 782 459 841 497
rect 782 425 788 459
rect 822 425 841 459
rect 782 387 841 425
rect 782 353 788 387
rect 822 353 841 387
rect 782 315 841 353
rect 782 281 788 315
rect 822 281 841 315
rect 782 243 841 281
rect 782 209 788 243
rect 822 209 841 243
rect 782 197 841 209
rect 264 125 618 137
rect 264 19 280 125
rect 602 19 618 125
rect 264 0 618 19
<< via1 >>
rect 203 603 255 639
rect 203 587 212 603
rect 212 587 246 603
rect 246 587 255 603
rect 203 569 212 575
rect 212 569 246 575
rect 246 569 255 575
rect 203 531 255 569
rect 203 523 212 531
rect 212 523 246 531
rect 246 523 255 531
rect 203 497 212 511
rect 212 497 246 511
rect 246 497 255 511
rect 203 459 255 497
rect 203 425 212 447
rect 212 425 246 447
rect 246 425 255 447
rect 203 395 255 425
rect 203 353 212 383
rect 212 353 246 383
rect 246 353 255 383
rect 203 331 255 353
rect 203 315 255 319
rect 203 281 212 315
rect 212 281 246 315
rect 246 281 255 315
rect 203 267 255 281
rect 203 243 255 255
rect 203 209 212 243
rect 212 209 246 243
rect 246 209 255 243
rect 203 203 255 209
rect 309 1179 361 1185
rect 309 1145 318 1179
rect 318 1145 352 1179
rect 352 1145 361 1179
rect 309 1133 361 1145
rect 309 1107 361 1121
rect 309 1073 318 1107
rect 318 1073 352 1107
rect 352 1073 361 1107
rect 309 1069 361 1073
rect 309 1035 361 1057
rect 309 1005 318 1035
rect 318 1005 352 1035
rect 352 1005 361 1035
rect 309 963 361 993
rect 309 941 318 963
rect 318 941 352 963
rect 352 941 361 963
rect 309 891 361 929
rect 309 877 318 891
rect 318 877 352 891
rect 352 877 361 891
rect 309 857 318 865
rect 318 857 352 865
rect 352 857 361 865
rect 309 819 361 857
rect 309 813 318 819
rect 318 813 352 819
rect 352 813 361 819
rect 309 785 318 801
rect 318 785 352 801
rect 352 785 361 801
rect 309 749 361 785
rect 415 603 467 639
rect 415 587 424 603
rect 424 587 458 603
rect 458 587 467 603
rect 415 569 424 575
rect 424 569 458 575
rect 458 569 467 575
rect 415 531 467 569
rect 415 523 424 531
rect 424 523 458 531
rect 458 523 467 531
rect 415 497 424 511
rect 424 497 458 511
rect 458 497 467 511
rect 415 459 467 497
rect 415 425 424 447
rect 424 425 458 447
rect 458 425 467 447
rect 415 395 467 425
rect 415 353 424 383
rect 424 353 458 383
rect 458 353 467 383
rect 415 331 467 353
rect 415 315 467 319
rect 415 281 424 315
rect 424 281 458 315
rect 458 281 467 315
rect 415 267 467 281
rect 415 243 467 255
rect 415 209 424 243
rect 424 209 458 243
rect 458 209 467 243
rect 415 203 467 209
rect 521 1179 573 1185
rect 521 1145 530 1179
rect 530 1145 564 1179
rect 564 1145 573 1179
rect 521 1133 573 1145
rect 521 1107 573 1121
rect 521 1073 530 1107
rect 530 1073 564 1107
rect 564 1073 573 1107
rect 521 1069 573 1073
rect 521 1035 573 1057
rect 521 1005 530 1035
rect 530 1005 564 1035
rect 564 1005 573 1035
rect 521 963 573 993
rect 521 941 530 963
rect 530 941 564 963
rect 564 941 573 963
rect 521 891 573 929
rect 521 877 530 891
rect 530 877 564 891
rect 564 877 573 891
rect 521 857 530 865
rect 530 857 564 865
rect 564 857 573 865
rect 521 819 573 857
rect 521 813 530 819
rect 530 813 564 819
rect 564 813 573 819
rect 521 785 530 801
rect 530 785 564 801
rect 564 785 573 801
rect 521 749 573 785
rect 627 603 679 639
rect 627 587 636 603
rect 636 587 670 603
rect 670 587 679 603
rect 627 569 636 575
rect 636 569 670 575
rect 670 569 679 575
rect 627 531 679 569
rect 627 523 636 531
rect 636 523 670 531
rect 670 523 679 531
rect 627 497 636 511
rect 636 497 670 511
rect 670 497 679 511
rect 627 459 679 497
rect 627 425 636 447
rect 636 425 670 447
rect 670 425 679 447
rect 627 395 679 425
rect 627 353 636 383
rect 636 353 670 383
rect 670 353 679 383
rect 627 331 679 353
rect 627 315 679 319
rect 627 281 636 315
rect 636 281 670 315
rect 670 281 679 315
rect 627 267 679 281
rect 627 243 679 255
rect 627 209 636 243
rect 636 209 670 243
rect 670 209 679 243
rect 627 203 679 209
<< metal2 >>
rect 14 1185 868 1191
rect 14 1133 309 1185
rect 361 1133 521 1185
rect 573 1133 868 1185
rect 14 1121 868 1133
rect 14 1069 309 1121
rect 361 1069 521 1121
rect 573 1069 868 1121
rect 14 1057 868 1069
rect 14 1005 309 1057
rect 361 1005 521 1057
rect 573 1005 868 1057
rect 14 993 868 1005
rect 14 941 309 993
rect 361 941 521 993
rect 573 941 868 993
rect 14 929 868 941
rect 14 877 309 929
rect 361 877 521 929
rect 573 877 868 929
rect 14 865 868 877
rect 14 813 309 865
rect 361 813 521 865
rect 573 813 868 865
rect 14 801 868 813
rect 14 749 309 801
rect 361 749 521 801
rect 573 749 868 801
rect 14 719 868 749
rect 14 639 868 669
rect 14 587 203 639
rect 255 587 415 639
rect 467 587 627 639
rect 679 587 868 639
rect 14 575 868 587
rect 14 523 203 575
rect 255 523 415 575
rect 467 523 627 575
rect 679 523 868 575
rect 14 511 868 523
rect 14 459 203 511
rect 255 459 415 511
rect 467 459 627 511
rect 679 459 868 511
rect 14 447 868 459
rect 14 395 203 447
rect 255 395 415 447
rect 467 395 627 447
rect 679 395 868 447
rect 14 383 868 395
rect 14 331 203 383
rect 255 331 415 383
rect 467 331 627 383
rect 679 331 868 383
rect 14 319 868 331
rect 14 267 203 319
rect 255 267 415 319
rect 467 267 627 319
rect 679 267 868 319
rect 14 255 868 267
rect 14 203 203 255
rect 255 203 415 255
rect 467 203 627 255
rect 679 203 868 255
rect 14 197 868 203
<< labels >>
flabel metal1 s 321 42 571 92 0 FreeSans 200 0 0 0 GATE
port 3 nsew
flabel metal1 s 321 1286 571 1336 0 FreeSans 200 0 0 0 GATE
port 3 nsew
flabel metal1 s 41 675 100 705 0 FreeSans 200 90 0 0 BULK
port 1 nsew
flabel metal1 s 782 683 841 713 0 FreeSans 200 90 0 0 BULK
port 1 nsew
flabel comment s 184 710 184 710 0 FreeSans 200 90 0 0 dummy_poly
flabel comment s 693 726 693 726 0 FreeSans 200 90 0 0 dummy_poly
flabel comment s 355 694 355 694 0 FreeSans 300 0 0 0 D
flabel comment s 269 694 269 694 0 FreeSans 300 0 0 0 S
flabel comment s 527 694 527 694 0 FreeSans 300 0 0 0 S
flabel comment s 441 694 441 694 0 FreeSans 300 0 0 0 S
flabel comment s 355 694 355 694 0 FreeSans 300 0 0 0 S
flabel comment s 269 694 269 694 0 FreeSans 300 0 0 0 S
flabel comment s 613 694 613 694 0 FreeSans 300 0 0 0 S
flabel comment s 527 694 527 694 0 FreeSans 300 0 0 0 D
flabel comment s 441 694 441 694 0 FreeSans 300 0 0 0 S
flabel metal2 s 14 384 35 512 7 FreeSans 300 180 0 0 SOURCE
port 4 nsew
flabel metal2 s 14 908 35 1036 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9880362
string GDS_START 9852188
<< end >>

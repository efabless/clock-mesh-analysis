magic
tech sky130A
magscale 1 2
timestamp 1633016076
<< checkpaint >>
rect -1260 -1260 3252 3852
<< dnwell >>
rect 214 214 1778 2378
<< nwell >>
rect 134 2098 1858 2458
rect 134 494 494 2098
rect 1498 494 1858 2098
rect 134 134 1858 494
<< pwell >>
rect 0 2458 1992 2592
rect 0 134 134 2458
rect 628 628 1364 1964
rect 1858 134 1992 2458
rect 0 0 1992 134
<< ndiff >>
rect 896 1653 1096 1696
rect 896 939 911 1653
rect 1081 939 1096 1653
rect 896 896 1096 939
<< ndiffc >>
rect 911 939 1081 1653
<< psubdiff >>
rect 26 2542 1966 2566
rect 26 2508 50 2542
rect 84 2508 129 2542
rect 163 2508 197 2542
rect 231 2508 265 2542
rect 299 2508 333 2542
rect 367 2508 401 2542
rect 435 2508 469 2542
rect 503 2508 537 2542
rect 571 2508 605 2542
rect 639 2508 673 2542
rect 707 2508 741 2542
rect 775 2508 809 2542
rect 843 2508 877 2542
rect 911 2508 945 2542
rect 979 2508 1013 2542
rect 1047 2508 1081 2542
rect 1115 2508 1149 2542
rect 1183 2508 1217 2542
rect 1251 2508 1285 2542
rect 1319 2508 1353 2542
rect 1387 2508 1421 2542
rect 1455 2508 1489 2542
rect 1523 2508 1557 2542
rect 1591 2508 1625 2542
rect 1659 2508 1693 2542
rect 1727 2508 1761 2542
rect 1795 2508 1829 2542
rect 1863 2508 1908 2542
rect 1942 2508 1966 2542
rect 26 2484 1966 2508
rect 26 2469 108 2484
rect 26 2435 50 2469
rect 84 2435 108 2469
rect 26 2401 108 2435
rect 26 2367 50 2401
rect 84 2367 108 2401
rect 26 2333 108 2367
rect 1884 2469 1966 2484
rect 1884 2435 1908 2469
rect 1942 2435 1966 2469
rect 1884 2401 1966 2435
rect 1884 2367 1908 2401
rect 1942 2367 1966 2401
rect 26 2299 50 2333
rect 84 2299 108 2333
rect 26 2265 108 2299
rect 26 2231 50 2265
rect 84 2231 108 2265
rect 26 2197 108 2231
rect 26 2163 50 2197
rect 84 2163 108 2197
rect 26 2129 108 2163
rect 26 2095 50 2129
rect 84 2095 108 2129
rect 26 2061 108 2095
rect 26 2027 50 2061
rect 84 2027 108 2061
rect 26 1993 108 2027
rect 26 1959 50 1993
rect 84 1959 108 1993
rect 26 1925 108 1959
rect 26 1891 50 1925
rect 84 1891 108 1925
rect 26 1857 108 1891
rect 26 1823 50 1857
rect 84 1823 108 1857
rect 26 1789 108 1823
rect 26 1755 50 1789
rect 84 1755 108 1789
rect 26 1721 108 1755
rect 26 1687 50 1721
rect 84 1687 108 1721
rect 26 1653 108 1687
rect 26 1619 50 1653
rect 84 1619 108 1653
rect 26 1585 108 1619
rect 26 1551 50 1585
rect 84 1551 108 1585
rect 26 1517 108 1551
rect 26 1483 50 1517
rect 84 1483 108 1517
rect 26 1449 108 1483
rect 26 1415 50 1449
rect 84 1415 108 1449
rect 26 1381 108 1415
rect 26 1347 50 1381
rect 84 1347 108 1381
rect 26 1313 108 1347
rect 26 1279 50 1313
rect 84 1279 108 1313
rect 26 1245 108 1279
rect 26 1211 50 1245
rect 84 1211 108 1245
rect 26 1177 108 1211
rect 26 1143 50 1177
rect 84 1143 108 1177
rect 26 1109 108 1143
rect 26 1075 50 1109
rect 84 1075 108 1109
rect 26 1041 108 1075
rect 26 1007 50 1041
rect 84 1007 108 1041
rect 26 973 108 1007
rect 26 939 50 973
rect 84 939 108 973
rect 26 905 108 939
rect 26 871 50 905
rect 84 871 108 905
rect 26 837 108 871
rect 26 803 50 837
rect 84 803 108 837
rect 26 769 108 803
rect 26 735 50 769
rect 84 735 108 769
rect 26 701 108 735
rect 26 667 50 701
rect 84 667 108 701
rect 26 633 108 667
rect 26 599 50 633
rect 84 599 108 633
rect 26 565 108 599
rect 26 531 50 565
rect 84 531 108 565
rect 26 497 108 531
rect 26 463 50 497
rect 84 463 108 497
rect 26 429 108 463
rect 26 395 50 429
rect 84 395 108 429
rect 26 361 108 395
rect 26 327 50 361
rect 84 327 108 361
rect 26 293 108 327
rect 26 259 50 293
rect 84 259 108 293
rect 26 225 108 259
rect 654 1914 1338 1938
rect 654 1880 678 1914
rect 712 1880 775 1914
rect 809 1880 843 1914
rect 877 1880 911 1914
rect 945 1880 979 1914
rect 1013 1880 1047 1914
rect 1081 1880 1115 1914
rect 1149 1880 1183 1914
rect 1217 1880 1280 1914
rect 1314 1880 1338 1914
rect 654 1856 1338 1880
rect 654 1823 736 1856
rect 654 1789 678 1823
rect 712 1789 736 1823
rect 654 1755 736 1789
rect 654 1721 678 1755
rect 712 1721 736 1755
rect 654 1687 736 1721
rect 1256 1823 1338 1856
rect 1256 1789 1280 1823
rect 1314 1789 1338 1823
rect 1256 1755 1338 1789
rect 1256 1721 1280 1755
rect 1314 1721 1338 1755
rect 654 1653 678 1687
rect 712 1653 736 1687
rect 654 1619 736 1653
rect 654 1585 678 1619
rect 712 1585 736 1619
rect 654 1551 736 1585
rect 654 1517 678 1551
rect 712 1517 736 1551
rect 654 1483 736 1517
rect 654 1449 678 1483
rect 712 1449 736 1483
rect 654 1415 736 1449
rect 654 1381 678 1415
rect 712 1381 736 1415
rect 654 1347 736 1381
rect 654 1313 678 1347
rect 712 1313 736 1347
rect 654 1279 736 1313
rect 654 1245 678 1279
rect 712 1245 736 1279
rect 654 1211 736 1245
rect 654 1177 678 1211
rect 712 1177 736 1211
rect 654 1143 736 1177
rect 654 1109 678 1143
rect 712 1109 736 1143
rect 654 1075 736 1109
rect 654 1041 678 1075
rect 712 1041 736 1075
rect 654 1007 736 1041
rect 654 973 678 1007
rect 712 973 736 1007
rect 654 939 736 973
rect 654 905 678 939
rect 712 905 736 939
rect 654 871 736 905
rect 1256 1687 1338 1721
rect 1256 1653 1280 1687
rect 1314 1653 1338 1687
rect 1256 1619 1338 1653
rect 1256 1585 1280 1619
rect 1314 1585 1338 1619
rect 1256 1551 1338 1585
rect 1256 1517 1280 1551
rect 1314 1517 1338 1551
rect 1256 1483 1338 1517
rect 1256 1449 1280 1483
rect 1314 1449 1338 1483
rect 1256 1415 1338 1449
rect 1256 1381 1280 1415
rect 1314 1381 1338 1415
rect 1256 1347 1338 1381
rect 1256 1313 1280 1347
rect 1314 1313 1338 1347
rect 1256 1279 1338 1313
rect 1256 1245 1280 1279
rect 1314 1245 1338 1279
rect 1256 1211 1338 1245
rect 1256 1177 1280 1211
rect 1314 1177 1338 1211
rect 1256 1143 1338 1177
rect 1256 1109 1280 1143
rect 1314 1109 1338 1143
rect 1256 1075 1338 1109
rect 1256 1041 1280 1075
rect 1314 1041 1338 1075
rect 1256 1007 1338 1041
rect 1256 973 1280 1007
rect 1314 973 1338 1007
rect 1256 939 1338 973
rect 1256 905 1280 939
rect 1314 905 1338 939
rect 654 837 678 871
rect 712 837 736 871
rect 654 803 736 837
rect 654 769 678 803
rect 712 769 736 803
rect 654 736 736 769
rect 1256 871 1338 905
rect 1256 837 1280 871
rect 1314 837 1338 871
rect 1256 803 1338 837
rect 1256 769 1280 803
rect 1314 769 1338 803
rect 1256 736 1338 769
rect 654 712 1338 736
rect 654 678 678 712
rect 712 678 775 712
rect 809 678 843 712
rect 877 678 911 712
rect 945 678 979 712
rect 1013 678 1047 712
rect 1081 678 1115 712
rect 1149 678 1183 712
rect 1217 678 1280 712
rect 1314 678 1338 712
rect 654 654 1338 678
rect 1884 2333 1966 2367
rect 1884 2299 1908 2333
rect 1942 2299 1966 2333
rect 1884 2265 1966 2299
rect 1884 2231 1908 2265
rect 1942 2231 1966 2265
rect 1884 2197 1966 2231
rect 1884 2163 1908 2197
rect 1942 2163 1966 2197
rect 1884 2129 1966 2163
rect 1884 2095 1908 2129
rect 1942 2095 1966 2129
rect 1884 2061 1966 2095
rect 1884 2027 1908 2061
rect 1942 2027 1966 2061
rect 1884 1993 1966 2027
rect 1884 1959 1908 1993
rect 1942 1959 1966 1993
rect 1884 1925 1966 1959
rect 1884 1891 1908 1925
rect 1942 1891 1966 1925
rect 1884 1857 1966 1891
rect 1884 1823 1908 1857
rect 1942 1823 1966 1857
rect 1884 1789 1966 1823
rect 1884 1755 1908 1789
rect 1942 1755 1966 1789
rect 1884 1721 1966 1755
rect 1884 1687 1908 1721
rect 1942 1687 1966 1721
rect 1884 1653 1966 1687
rect 1884 1619 1908 1653
rect 1942 1619 1966 1653
rect 1884 1585 1966 1619
rect 1884 1551 1908 1585
rect 1942 1551 1966 1585
rect 1884 1517 1966 1551
rect 1884 1483 1908 1517
rect 1942 1483 1966 1517
rect 1884 1449 1966 1483
rect 1884 1415 1908 1449
rect 1942 1415 1966 1449
rect 1884 1381 1966 1415
rect 1884 1347 1908 1381
rect 1942 1347 1966 1381
rect 1884 1313 1966 1347
rect 1884 1279 1908 1313
rect 1942 1279 1966 1313
rect 1884 1245 1966 1279
rect 1884 1211 1908 1245
rect 1942 1211 1966 1245
rect 1884 1177 1966 1211
rect 1884 1143 1908 1177
rect 1942 1143 1966 1177
rect 1884 1109 1966 1143
rect 1884 1075 1908 1109
rect 1942 1075 1966 1109
rect 1884 1041 1966 1075
rect 1884 1007 1908 1041
rect 1942 1007 1966 1041
rect 1884 973 1966 1007
rect 1884 939 1908 973
rect 1942 939 1966 973
rect 1884 905 1966 939
rect 1884 871 1908 905
rect 1942 871 1966 905
rect 1884 837 1966 871
rect 1884 803 1908 837
rect 1942 803 1966 837
rect 1884 769 1966 803
rect 1884 735 1908 769
rect 1942 735 1966 769
rect 1884 701 1966 735
rect 1884 667 1908 701
rect 1942 667 1966 701
rect 1884 633 1966 667
rect 1884 599 1908 633
rect 1942 599 1966 633
rect 1884 565 1966 599
rect 1884 531 1908 565
rect 1942 531 1966 565
rect 1884 497 1966 531
rect 1884 463 1908 497
rect 1942 463 1966 497
rect 1884 429 1966 463
rect 1884 395 1908 429
rect 1942 395 1966 429
rect 1884 361 1966 395
rect 1884 327 1908 361
rect 1942 327 1966 361
rect 1884 293 1966 327
rect 1884 259 1908 293
rect 1942 259 1966 293
rect 26 191 50 225
rect 84 191 108 225
rect 26 157 108 191
rect 26 123 50 157
rect 84 123 108 157
rect 26 108 108 123
rect 1884 225 1966 259
rect 1884 191 1908 225
rect 1942 191 1966 225
rect 1884 157 1966 191
rect 1884 123 1908 157
rect 1942 123 1966 157
rect 1884 108 1966 123
rect 26 84 1966 108
rect 26 50 50 84
rect 84 50 129 84
rect 163 50 197 84
rect 231 50 265 84
rect 299 50 333 84
rect 367 50 401 84
rect 435 50 469 84
rect 503 50 537 84
rect 571 50 605 84
rect 639 50 673 84
rect 707 50 741 84
rect 775 50 809 84
rect 843 50 877 84
rect 911 50 945 84
rect 979 50 1013 84
rect 1047 50 1081 84
rect 1115 50 1149 84
rect 1183 50 1217 84
rect 1251 50 1285 84
rect 1319 50 1353 84
rect 1387 50 1421 84
rect 1455 50 1489 84
rect 1523 50 1557 84
rect 1591 50 1625 84
rect 1659 50 1693 84
rect 1727 50 1761 84
rect 1795 50 1829 84
rect 1863 50 1908 84
rect 1942 50 1966 84
rect 26 26 1966 50
<< nsubdiff >>
rect 252 2316 1740 2340
rect 252 2282 276 2316
rect 310 2282 367 2316
rect 401 2282 435 2316
rect 469 2282 503 2316
rect 537 2282 571 2316
rect 605 2282 639 2316
rect 673 2282 707 2316
rect 741 2282 775 2316
rect 809 2282 843 2316
rect 877 2282 911 2316
rect 945 2282 979 2316
rect 1013 2282 1047 2316
rect 1081 2282 1115 2316
rect 1149 2282 1183 2316
rect 1217 2282 1251 2316
rect 1285 2282 1319 2316
rect 1353 2282 1387 2316
rect 1421 2282 1455 2316
rect 1489 2282 1523 2316
rect 1557 2282 1591 2316
rect 1625 2282 1682 2316
rect 1716 2282 1740 2316
rect 252 2258 1740 2282
rect 252 2231 334 2258
rect 252 2197 276 2231
rect 310 2197 334 2231
rect 252 2163 334 2197
rect 252 2129 276 2163
rect 310 2129 334 2163
rect 252 2095 334 2129
rect 252 2061 276 2095
rect 310 2061 334 2095
rect 252 2027 334 2061
rect 252 1993 276 2027
rect 310 1993 334 2027
rect 252 1959 334 1993
rect 252 1925 276 1959
rect 310 1925 334 1959
rect 1658 2231 1740 2258
rect 1658 2197 1682 2231
rect 1716 2197 1740 2231
rect 1658 2163 1740 2197
rect 1658 2129 1682 2163
rect 1716 2129 1740 2163
rect 1658 2095 1740 2129
rect 1658 2061 1682 2095
rect 1716 2061 1740 2095
rect 1658 2027 1740 2061
rect 1658 1993 1682 2027
rect 1716 1993 1740 2027
rect 1658 1959 1740 1993
rect 252 1891 334 1925
rect 252 1857 276 1891
rect 310 1857 334 1891
rect 252 1823 334 1857
rect 252 1789 276 1823
rect 310 1789 334 1823
rect 252 1755 334 1789
rect 252 1721 276 1755
rect 310 1721 334 1755
rect 252 1687 334 1721
rect 252 1653 276 1687
rect 310 1653 334 1687
rect 252 1619 334 1653
rect 252 1585 276 1619
rect 310 1585 334 1619
rect 252 1551 334 1585
rect 252 1517 276 1551
rect 310 1517 334 1551
rect 252 1483 334 1517
rect 252 1449 276 1483
rect 310 1449 334 1483
rect 252 1415 334 1449
rect 252 1381 276 1415
rect 310 1381 334 1415
rect 252 1347 334 1381
rect 252 1313 276 1347
rect 310 1313 334 1347
rect 252 1279 334 1313
rect 252 1245 276 1279
rect 310 1245 334 1279
rect 252 1211 334 1245
rect 252 1177 276 1211
rect 310 1177 334 1211
rect 252 1143 334 1177
rect 252 1109 276 1143
rect 310 1109 334 1143
rect 252 1075 334 1109
rect 252 1041 276 1075
rect 310 1041 334 1075
rect 252 1007 334 1041
rect 252 973 276 1007
rect 310 973 334 1007
rect 252 939 334 973
rect 252 905 276 939
rect 310 905 334 939
rect 252 871 334 905
rect 252 837 276 871
rect 310 837 334 871
rect 252 803 334 837
rect 252 769 276 803
rect 310 769 334 803
rect 252 735 334 769
rect 252 701 276 735
rect 310 701 334 735
rect 252 667 334 701
rect 252 633 276 667
rect 310 633 334 667
rect 1658 1925 1682 1959
rect 1716 1925 1740 1959
rect 1658 1891 1740 1925
rect 1658 1857 1682 1891
rect 1716 1857 1740 1891
rect 1658 1823 1740 1857
rect 1658 1789 1682 1823
rect 1716 1789 1740 1823
rect 1658 1755 1740 1789
rect 1658 1721 1682 1755
rect 1716 1721 1740 1755
rect 1658 1687 1740 1721
rect 1658 1653 1682 1687
rect 1716 1653 1740 1687
rect 1658 1619 1740 1653
rect 1658 1585 1682 1619
rect 1716 1585 1740 1619
rect 1658 1551 1740 1585
rect 1658 1517 1682 1551
rect 1716 1517 1740 1551
rect 1658 1483 1740 1517
rect 1658 1449 1682 1483
rect 1716 1449 1740 1483
rect 1658 1415 1740 1449
rect 1658 1381 1682 1415
rect 1716 1381 1740 1415
rect 1658 1347 1740 1381
rect 1658 1313 1682 1347
rect 1716 1313 1740 1347
rect 1658 1279 1740 1313
rect 1658 1245 1682 1279
rect 1716 1245 1740 1279
rect 1658 1211 1740 1245
rect 1658 1177 1682 1211
rect 1716 1177 1740 1211
rect 1658 1143 1740 1177
rect 1658 1109 1682 1143
rect 1716 1109 1740 1143
rect 1658 1075 1740 1109
rect 1658 1041 1682 1075
rect 1716 1041 1740 1075
rect 1658 1007 1740 1041
rect 1658 973 1682 1007
rect 1716 973 1740 1007
rect 1658 939 1740 973
rect 1658 905 1682 939
rect 1716 905 1740 939
rect 1658 871 1740 905
rect 1658 837 1682 871
rect 1716 837 1740 871
rect 1658 803 1740 837
rect 1658 769 1682 803
rect 1716 769 1740 803
rect 1658 735 1740 769
rect 1658 701 1682 735
rect 1716 701 1740 735
rect 1658 667 1740 701
rect 252 599 334 633
rect 252 565 276 599
rect 310 565 334 599
rect 252 531 334 565
rect 252 497 276 531
rect 310 497 334 531
rect 252 463 334 497
rect 252 429 276 463
rect 310 429 334 463
rect 252 395 334 429
rect 252 361 276 395
rect 310 361 334 395
rect 252 334 334 361
rect 1658 633 1682 667
rect 1716 633 1740 667
rect 1658 599 1740 633
rect 1658 565 1682 599
rect 1716 565 1740 599
rect 1658 531 1740 565
rect 1658 497 1682 531
rect 1716 497 1740 531
rect 1658 463 1740 497
rect 1658 429 1682 463
rect 1716 429 1740 463
rect 1658 395 1740 429
rect 1658 361 1682 395
rect 1716 361 1740 395
rect 1658 334 1740 361
rect 252 310 1740 334
rect 252 276 276 310
rect 310 276 367 310
rect 401 276 435 310
rect 469 276 503 310
rect 537 276 571 310
rect 605 276 639 310
rect 673 276 707 310
rect 741 276 775 310
rect 809 276 843 310
rect 877 276 911 310
rect 945 276 979 310
rect 1013 276 1047 310
rect 1081 276 1115 310
rect 1149 276 1183 310
rect 1217 276 1251 310
rect 1285 276 1319 310
rect 1353 276 1387 310
rect 1421 276 1455 310
rect 1489 276 1523 310
rect 1557 276 1591 310
rect 1625 276 1682 310
rect 1716 276 1740 310
rect 252 252 1740 276
<< psubdiffcont >>
rect 50 2508 84 2542
rect 129 2508 163 2542
rect 197 2508 231 2542
rect 265 2508 299 2542
rect 333 2508 367 2542
rect 401 2508 435 2542
rect 469 2508 503 2542
rect 537 2508 571 2542
rect 605 2508 639 2542
rect 673 2508 707 2542
rect 741 2508 775 2542
rect 809 2508 843 2542
rect 877 2508 911 2542
rect 945 2508 979 2542
rect 1013 2508 1047 2542
rect 1081 2508 1115 2542
rect 1149 2508 1183 2542
rect 1217 2508 1251 2542
rect 1285 2508 1319 2542
rect 1353 2508 1387 2542
rect 1421 2508 1455 2542
rect 1489 2508 1523 2542
rect 1557 2508 1591 2542
rect 1625 2508 1659 2542
rect 1693 2508 1727 2542
rect 1761 2508 1795 2542
rect 1829 2508 1863 2542
rect 1908 2508 1942 2542
rect 50 2435 84 2469
rect 50 2367 84 2401
rect 1908 2435 1942 2469
rect 1908 2367 1942 2401
rect 50 2299 84 2333
rect 50 2231 84 2265
rect 50 2163 84 2197
rect 50 2095 84 2129
rect 50 2027 84 2061
rect 50 1959 84 1993
rect 50 1891 84 1925
rect 50 1823 84 1857
rect 50 1755 84 1789
rect 50 1687 84 1721
rect 50 1619 84 1653
rect 50 1551 84 1585
rect 50 1483 84 1517
rect 50 1415 84 1449
rect 50 1347 84 1381
rect 50 1279 84 1313
rect 50 1211 84 1245
rect 50 1143 84 1177
rect 50 1075 84 1109
rect 50 1007 84 1041
rect 50 939 84 973
rect 50 871 84 905
rect 50 803 84 837
rect 50 735 84 769
rect 50 667 84 701
rect 50 599 84 633
rect 50 531 84 565
rect 50 463 84 497
rect 50 395 84 429
rect 50 327 84 361
rect 50 259 84 293
rect 678 1880 712 1914
rect 775 1880 809 1914
rect 843 1880 877 1914
rect 911 1880 945 1914
rect 979 1880 1013 1914
rect 1047 1880 1081 1914
rect 1115 1880 1149 1914
rect 1183 1880 1217 1914
rect 1280 1880 1314 1914
rect 678 1789 712 1823
rect 678 1721 712 1755
rect 1280 1789 1314 1823
rect 1280 1721 1314 1755
rect 678 1653 712 1687
rect 678 1585 712 1619
rect 678 1517 712 1551
rect 678 1449 712 1483
rect 678 1381 712 1415
rect 678 1313 712 1347
rect 678 1245 712 1279
rect 678 1177 712 1211
rect 678 1109 712 1143
rect 678 1041 712 1075
rect 678 973 712 1007
rect 678 905 712 939
rect 1280 1653 1314 1687
rect 1280 1585 1314 1619
rect 1280 1517 1314 1551
rect 1280 1449 1314 1483
rect 1280 1381 1314 1415
rect 1280 1313 1314 1347
rect 1280 1245 1314 1279
rect 1280 1177 1314 1211
rect 1280 1109 1314 1143
rect 1280 1041 1314 1075
rect 1280 973 1314 1007
rect 1280 905 1314 939
rect 678 837 712 871
rect 678 769 712 803
rect 1280 837 1314 871
rect 1280 769 1314 803
rect 678 678 712 712
rect 775 678 809 712
rect 843 678 877 712
rect 911 678 945 712
rect 979 678 1013 712
rect 1047 678 1081 712
rect 1115 678 1149 712
rect 1183 678 1217 712
rect 1280 678 1314 712
rect 1908 2299 1942 2333
rect 1908 2231 1942 2265
rect 1908 2163 1942 2197
rect 1908 2095 1942 2129
rect 1908 2027 1942 2061
rect 1908 1959 1942 1993
rect 1908 1891 1942 1925
rect 1908 1823 1942 1857
rect 1908 1755 1942 1789
rect 1908 1687 1942 1721
rect 1908 1619 1942 1653
rect 1908 1551 1942 1585
rect 1908 1483 1942 1517
rect 1908 1415 1942 1449
rect 1908 1347 1942 1381
rect 1908 1279 1942 1313
rect 1908 1211 1942 1245
rect 1908 1143 1942 1177
rect 1908 1075 1942 1109
rect 1908 1007 1942 1041
rect 1908 939 1942 973
rect 1908 871 1942 905
rect 1908 803 1942 837
rect 1908 735 1942 769
rect 1908 667 1942 701
rect 1908 599 1942 633
rect 1908 531 1942 565
rect 1908 463 1942 497
rect 1908 395 1942 429
rect 1908 327 1942 361
rect 1908 259 1942 293
rect 50 191 84 225
rect 50 123 84 157
rect 1908 191 1942 225
rect 1908 123 1942 157
rect 50 50 84 84
rect 129 50 163 84
rect 197 50 231 84
rect 265 50 299 84
rect 333 50 367 84
rect 401 50 435 84
rect 469 50 503 84
rect 537 50 571 84
rect 605 50 639 84
rect 673 50 707 84
rect 741 50 775 84
rect 809 50 843 84
rect 877 50 911 84
rect 945 50 979 84
rect 1013 50 1047 84
rect 1081 50 1115 84
rect 1149 50 1183 84
rect 1217 50 1251 84
rect 1285 50 1319 84
rect 1353 50 1387 84
rect 1421 50 1455 84
rect 1489 50 1523 84
rect 1557 50 1591 84
rect 1625 50 1659 84
rect 1693 50 1727 84
rect 1761 50 1795 84
rect 1829 50 1863 84
rect 1908 50 1942 84
<< nsubdiffcont >>
rect 276 2282 310 2316
rect 367 2282 401 2316
rect 435 2282 469 2316
rect 503 2282 537 2316
rect 571 2282 605 2316
rect 639 2282 673 2316
rect 707 2282 741 2316
rect 775 2282 809 2316
rect 843 2282 877 2316
rect 911 2282 945 2316
rect 979 2282 1013 2316
rect 1047 2282 1081 2316
rect 1115 2282 1149 2316
rect 1183 2282 1217 2316
rect 1251 2282 1285 2316
rect 1319 2282 1353 2316
rect 1387 2282 1421 2316
rect 1455 2282 1489 2316
rect 1523 2282 1557 2316
rect 1591 2282 1625 2316
rect 1682 2282 1716 2316
rect 276 2197 310 2231
rect 276 2129 310 2163
rect 276 2061 310 2095
rect 276 1993 310 2027
rect 276 1925 310 1959
rect 1682 2197 1716 2231
rect 1682 2129 1716 2163
rect 1682 2061 1716 2095
rect 1682 1993 1716 2027
rect 276 1857 310 1891
rect 276 1789 310 1823
rect 276 1721 310 1755
rect 276 1653 310 1687
rect 276 1585 310 1619
rect 276 1517 310 1551
rect 276 1449 310 1483
rect 276 1381 310 1415
rect 276 1313 310 1347
rect 276 1245 310 1279
rect 276 1177 310 1211
rect 276 1109 310 1143
rect 276 1041 310 1075
rect 276 973 310 1007
rect 276 905 310 939
rect 276 837 310 871
rect 276 769 310 803
rect 276 701 310 735
rect 276 633 310 667
rect 1682 1925 1716 1959
rect 1682 1857 1716 1891
rect 1682 1789 1716 1823
rect 1682 1721 1716 1755
rect 1682 1653 1716 1687
rect 1682 1585 1716 1619
rect 1682 1517 1716 1551
rect 1682 1449 1716 1483
rect 1682 1381 1716 1415
rect 1682 1313 1716 1347
rect 1682 1245 1716 1279
rect 1682 1177 1716 1211
rect 1682 1109 1716 1143
rect 1682 1041 1716 1075
rect 1682 973 1716 1007
rect 1682 905 1716 939
rect 1682 837 1716 871
rect 1682 769 1716 803
rect 1682 701 1716 735
rect 276 565 310 599
rect 276 497 310 531
rect 276 429 310 463
rect 276 361 310 395
rect 1682 633 1716 667
rect 1682 565 1716 599
rect 1682 497 1716 531
rect 1682 429 1716 463
rect 1682 361 1716 395
rect 276 276 310 310
rect 367 276 401 310
rect 435 276 469 310
rect 503 276 537 310
rect 571 276 605 310
rect 639 276 673 310
rect 707 276 741 310
rect 775 276 809 310
rect 843 276 877 310
rect 911 276 945 310
rect 979 276 1013 310
rect 1047 276 1081 310
rect 1115 276 1149 310
rect 1183 276 1217 310
rect 1251 276 1285 310
rect 1319 276 1353 310
rect 1387 276 1421 310
rect 1455 276 1489 310
rect 1523 276 1557 310
rect 1591 276 1625 310
rect 1682 276 1716 310
<< locali >>
rect 34 2542 1958 2558
rect 34 2508 50 2542
rect 84 2508 129 2542
rect 185 2508 197 2542
rect 257 2508 265 2542
rect 329 2508 333 2542
rect 435 2508 439 2542
rect 503 2508 511 2542
rect 571 2508 583 2542
rect 639 2508 655 2542
rect 707 2508 727 2542
rect 775 2508 799 2542
rect 843 2508 871 2542
rect 911 2508 943 2542
rect 979 2508 1013 2542
rect 1049 2508 1081 2542
rect 1121 2508 1149 2542
rect 1193 2508 1217 2542
rect 1265 2508 1285 2542
rect 1337 2508 1353 2542
rect 1409 2508 1421 2542
rect 1481 2508 1489 2542
rect 1553 2508 1557 2542
rect 1659 2508 1663 2542
rect 1727 2508 1735 2542
rect 1795 2508 1807 2542
rect 1863 2508 1908 2542
rect 1942 2508 1958 2542
rect 34 2492 1958 2508
rect 34 2469 100 2492
rect 34 2431 50 2469
rect 84 2431 100 2469
rect 34 2401 100 2431
rect 34 2359 50 2401
rect 84 2359 100 2401
rect 34 2333 100 2359
rect 34 2287 50 2333
rect 84 2287 100 2333
rect 1892 2469 1958 2492
rect 1892 2431 1908 2469
rect 1942 2431 1958 2469
rect 1892 2401 1958 2431
rect 1892 2359 1908 2401
rect 1942 2359 1958 2401
rect 1892 2333 1958 2359
rect 34 2265 100 2287
rect 34 2215 50 2265
rect 84 2215 100 2265
rect 34 2197 100 2215
rect 34 2143 50 2197
rect 84 2143 100 2197
rect 34 2129 100 2143
rect 34 2071 50 2129
rect 84 2071 100 2129
rect 34 2061 100 2071
rect 34 1999 50 2061
rect 84 1999 100 2061
rect 34 1993 100 1999
rect 34 1927 50 1993
rect 84 1927 100 1993
rect 34 1925 100 1927
rect 34 1891 50 1925
rect 84 1891 100 1925
rect 34 1889 100 1891
rect 34 1823 50 1889
rect 84 1823 100 1889
rect 34 1817 100 1823
rect 34 1755 50 1817
rect 84 1755 100 1817
rect 34 1745 100 1755
rect 34 1687 50 1745
rect 84 1687 100 1745
rect 34 1673 100 1687
rect 34 1619 50 1673
rect 84 1619 100 1673
rect 34 1601 100 1619
rect 34 1551 50 1601
rect 84 1551 100 1601
rect 34 1529 100 1551
rect 34 1483 50 1529
rect 84 1483 100 1529
rect 34 1457 100 1483
rect 34 1415 50 1457
rect 84 1415 100 1457
rect 34 1385 100 1415
rect 34 1347 50 1385
rect 84 1347 100 1385
rect 34 1313 100 1347
rect 34 1279 50 1313
rect 84 1279 100 1313
rect 34 1245 100 1279
rect 34 1207 50 1245
rect 84 1207 100 1245
rect 34 1177 100 1207
rect 34 1135 50 1177
rect 84 1135 100 1177
rect 34 1109 100 1135
rect 34 1063 50 1109
rect 84 1063 100 1109
rect 34 1041 100 1063
rect 34 991 50 1041
rect 84 991 100 1041
rect 34 973 100 991
rect 34 919 50 973
rect 84 919 100 973
rect 34 905 100 919
rect 34 847 50 905
rect 84 847 100 905
rect 34 837 100 847
rect 34 775 50 837
rect 84 775 100 837
rect 34 769 100 775
rect 34 703 50 769
rect 84 703 100 769
rect 34 701 100 703
rect 34 667 50 701
rect 84 667 100 701
rect 34 665 100 667
rect 34 599 50 665
rect 84 599 100 665
rect 34 593 100 599
rect 34 531 50 593
rect 84 531 100 593
rect 34 521 100 531
rect 34 463 50 521
rect 84 463 100 521
rect 34 449 100 463
rect 34 395 50 449
rect 84 395 100 449
rect 34 377 100 395
rect 34 327 50 377
rect 84 327 100 377
rect 34 305 100 327
rect 34 259 50 305
rect 84 259 100 305
rect 260 2316 1732 2332
rect 260 2282 276 2316
rect 310 2282 367 2316
rect 401 2282 435 2316
rect 473 2282 503 2316
rect 545 2282 571 2316
rect 617 2282 639 2316
rect 689 2282 707 2316
rect 761 2282 775 2316
rect 833 2282 843 2316
rect 905 2282 911 2316
rect 977 2282 979 2316
rect 1013 2282 1015 2316
rect 1081 2282 1087 2316
rect 1149 2282 1159 2316
rect 1217 2282 1231 2316
rect 1285 2282 1303 2316
rect 1353 2282 1375 2316
rect 1421 2282 1447 2316
rect 1489 2282 1519 2316
rect 1557 2282 1591 2316
rect 1625 2282 1682 2316
rect 1716 2282 1732 2316
rect 260 2266 1732 2282
rect 260 2231 326 2266
rect 260 2179 276 2231
rect 310 2179 326 2231
rect 260 2163 326 2179
rect 260 2107 276 2163
rect 310 2107 326 2163
rect 260 2095 326 2107
rect 260 2035 276 2095
rect 310 2035 326 2095
rect 260 2027 326 2035
rect 260 1963 276 2027
rect 310 1963 326 2027
rect 260 1959 326 1963
rect 260 1857 276 1959
rect 310 1857 326 1959
rect 1666 2231 1732 2266
rect 1666 2179 1682 2231
rect 1716 2179 1732 2231
rect 1666 2163 1732 2179
rect 1666 2107 1682 2163
rect 1716 2107 1732 2163
rect 1666 2095 1732 2107
rect 1666 2035 1682 2095
rect 1716 2035 1732 2095
rect 1666 2027 1732 2035
rect 1666 1963 1682 2027
rect 1716 1963 1732 2027
rect 1666 1959 1732 1963
rect 260 1853 326 1857
rect 260 1789 276 1853
rect 310 1789 326 1853
rect 260 1781 326 1789
rect 260 1721 276 1781
rect 310 1721 326 1781
rect 260 1709 326 1721
rect 260 1653 276 1709
rect 310 1653 326 1709
rect 260 1637 326 1653
rect 260 1585 276 1637
rect 310 1585 326 1637
rect 260 1565 326 1585
rect 260 1517 276 1565
rect 310 1517 326 1565
rect 260 1493 326 1517
rect 260 1449 276 1493
rect 310 1449 326 1493
rect 260 1421 326 1449
rect 260 1381 276 1421
rect 310 1381 326 1421
rect 260 1349 326 1381
rect 260 1313 276 1349
rect 310 1313 326 1349
rect 260 1279 326 1313
rect 260 1243 276 1279
rect 310 1243 326 1279
rect 260 1211 326 1243
rect 260 1171 276 1211
rect 310 1171 326 1211
rect 260 1143 326 1171
rect 260 1099 276 1143
rect 310 1099 326 1143
rect 260 1075 326 1099
rect 260 1027 276 1075
rect 310 1027 326 1075
rect 260 1007 326 1027
rect 260 955 276 1007
rect 310 955 326 1007
rect 260 939 326 955
rect 260 883 276 939
rect 310 883 326 939
rect 260 871 326 883
rect 260 811 276 871
rect 310 811 326 871
rect 260 803 326 811
rect 260 739 276 803
rect 310 739 326 803
rect 260 735 326 739
rect 260 633 276 735
rect 310 633 326 735
rect 662 1914 1330 1930
rect 662 1880 678 1914
rect 712 1880 763 1914
rect 809 1880 835 1914
rect 877 1880 907 1914
rect 945 1880 979 1914
rect 1013 1880 1047 1914
rect 1085 1880 1115 1914
rect 1157 1880 1183 1914
rect 1229 1880 1280 1914
rect 1314 1880 1330 1914
rect 662 1864 1330 1880
rect 662 1823 728 1864
rect 662 1783 678 1823
rect 712 1783 728 1823
rect 662 1755 728 1783
rect 662 1711 678 1755
rect 712 1711 728 1755
rect 662 1687 728 1711
rect 1264 1823 1330 1864
rect 1264 1783 1280 1823
rect 1314 1783 1330 1823
rect 1264 1755 1330 1783
rect 1264 1711 1280 1755
rect 1314 1711 1330 1755
rect 662 1639 678 1687
rect 712 1639 728 1687
rect 662 1619 728 1639
rect 662 1567 678 1619
rect 712 1567 728 1619
rect 662 1551 728 1567
rect 662 1495 678 1551
rect 712 1495 728 1551
rect 662 1483 728 1495
rect 662 1423 678 1483
rect 712 1423 728 1483
rect 662 1415 728 1423
rect 662 1351 678 1415
rect 712 1351 728 1415
rect 662 1347 728 1351
rect 662 1245 678 1347
rect 712 1245 728 1347
rect 662 1241 728 1245
rect 662 1177 678 1241
rect 712 1177 728 1241
rect 662 1169 728 1177
rect 662 1109 678 1169
rect 712 1109 728 1169
rect 662 1097 728 1109
rect 662 1041 678 1097
rect 712 1041 728 1097
rect 662 1025 728 1041
rect 662 973 678 1025
rect 712 973 728 1025
rect 662 953 728 973
rect 662 905 678 953
rect 712 905 728 953
rect 662 881 728 905
rect 895 1673 1097 1697
rect 895 919 907 1673
rect 1085 919 1097 1673
rect 895 895 1097 919
rect 1264 1687 1330 1711
rect 1264 1639 1280 1687
rect 1314 1639 1330 1687
rect 1264 1619 1330 1639
rect 1264 1567 1280 1619
rect 1314 1567 1330 1619
rect 1264 1551 1330 1567
rect 1264 1495 1280 1551
rect 1314 1495 1330 1551
rect 1264 1483 1330 1495
rect 1264 1423 1280 1483
rect 1314 1423 1330 1483
rect 1264 1415 1330 1423
rect 1264 1351 1280 1415
rect 1314 1351 1330 1415
rect 1264 1347 1330 1351
rect 1264 1245 1280 1347
rect 1314 1245 1330 1347
rect 1264 1241 1330 1245
rect 1264 1177 1280 1241
rect 1314 1177 1330 1241
rect 1264 1169 1330 1177
rect 1264 1109 1280 1169
rect 1314 1109 1330 1169
rect 1264 1097 1330 1109
rect 1264 1041 1280 1097
rect 1314 1041 1330 1097
rect 1264 1025 1330 1041
rect 1264 973 1280 1025
rect 1314 973 1330 1025
rect 1264 953 1330 973
rect 1264 905 1280 953
rect 1314 905 1330 953
rect 662 837 678 881
rect 712 837 728 881
rect 662 809 728 837
rect 662 769 678 809
rect 712 769 728 809
rect 662 728 728 769
rect 1264 881 1330 905
rect 1264 837 1280 881
rect 1314 837 1330 881
rect 1264 809 1330 837
rect 1264 769 1280 809
rect 1314 769 1330 809
rect 1264 728 1330 769
rect 662 712 1330 728
rect 662 678 678 712
rect 712 678 763 712
rect 809 678 835 712
rect 877 678 907 712
rect 945 678 979 712
rect 1013 678 1047 712
rect 1085 678 1115 712
rect 1157 678 1183 712
rect 1229 678 1280 712
rect 1314 678 1330 712
rect 662 662 1330 678
rect 1666 1857 1682 1959
rect 1716 1857 1732 1959
rect 1666 1853 1732 1857
rect 1666 1789 1682 1853
rect 1716 1789 1732 1853
rect 1666 1781 1732 1789
rect 1666 1721 1682 1781
rect 1716 1721 1732 1781
rect 1666 1709 1732 1721
rect 1666 1653 1682 1709
rect 1716 1653 1732 1709
rect 1666 1637 1732 1653
rect 1666 1585 1682 1637
rect 1716 1585 1732 1637
rect 1666 1565 1732 1585
rect 1666 1517 1682 1565
rect 1716 1517 1732 1565
rect 1666 1493 1732 1517
rect 1666 1449 1682 1493
rect 1716 1449 1732 1493
rect 1666 1421 1732 1449
rect 1666 1381 1682 1421
rect 1716 1381 1732 1421
rect 1666 1349 1732 1381
rect 1666 1313 1682 1349
rect 1716 1313 1732 1349
rect 1666 1279 1732 1313
rect 1666 1243 1682 1279
rect 1716 1243 1732 1279
rect 1666 1211 1732 1243
rect 1666 1171 1682 1211
rect 1716 1171 1732 1211
rect 1666 1143 1732 1171
rect 1666 1099 1682 1143
rect 1716 1099 1732 1143
rect 1666 1075 1732 1099
rect 1666 1027 1682 1075
rect 1716 1027 1732 1075
rect 1666 1007 1732 1027
rect 1666 955 1682 1007
rect 1716 955 1732 1007
rect 1666 939 1732 955
rect 1666 883 1682 939
rect 1716 883 1732 939
rect 1666 871 1732 883
rect 1666 811 1682 871
rect 1716 811 1732 871
rect 1666 803 1732 811
rect 1666 739 1682 803
rect 1716 739 1732 803
rect 1666 735 1732 739
rect 260 629 326 633
rect 260 565 276 629
rect 310 565 326 629
rect 260 557 326 565
rect 260 497 276 557
rect 310 497 326 557
rect 260 485 326 497
rect 260 429 276 485
rect 310 429 326 485
rect 260 413 326 429
rect 260 361 276 413
rect 310 361 326 413
rect 260 326 326 361
rect 1666 633 1682 735
rect 1716 633 1732 735
rect 1666 629 1732 633
rect 1666 565 1682 629
rect 1716 565 1732 629
rect 1666 557 1732 565
rect 1666 497 1682 557
rect 1716 497 1732 557
rect 1666 485 1732 497
rect 1666 429 1682 485
rect 1716 429 1732 485
rect 1666 413 1732 429
rect 1666 361 1682 413
rect 1716 361 1732 413
rect 1666 326 1732 361
rect 260 310 1732 326
rect 260 276 276 310
rect 310 276 367 310
rect 401 276 435 310
rect 473 276 503 310
rect 545 276 571 310
rect 617 276 639 310
rect 689 276 707 310
rect 761 276 775 310
rect 833 276 843 310
rect 905 276 911 310
rect 977 276 979 310
rect 1013 276 1015 310
rect 1081 276 1087 310
rect 1149 276 1159 310
rect 1217 276 1231 310
rect 1285 276 1303 310
rect 1353 276 1375 310
rect 1421 276 1447 310
rect 1489 276 1519 310
rect 1557 276 1591 310
rect 1625 276 1682 310
rect 1716 276 1732 310
rect 260 260 1732 276
rect 1892 2287 1908 2333
rect 1942 2287 1958 2333
rect 1892 2265 1958 2287
rect 1892 2215 1908 2265
rect 1942 2215 1958 2265
rect 1892 2197 1958 2215
rect 1892 2143 1908 2197
rect 1942 2143 1958 2197
rect 1892 2129 1958 2143
rect 1892 2071 1908 2129
rect 1942 2071 1958 2129
rect 1892 2061 1958 2071
rect 1892 1999 1908 2061
rect 1942 1999 1958 2061
rect 1892 1993 1958 1999
rect 1892 1927 1908 1993
rect 1942 1927 1958 1993
rect 1892 1925 1958 1927
rect 1892 1891 1908 1925
rect 1942 1891 1958 1925
rect 1892 1889 1958 1891
rect 1892 1823 1908 1889
rect 1942 1823 1958 1889
rect 1892 1817 1958 1823
rect 1892 1755 1908 1817
rect 1942 1755 1958 1817
rect 1892 1745 1958 1755
rect 1892 1687 1908 1745
rect 1942 1687 1958 1745
rect 1892 1673 1958 1687
rect 1892 1619 1908 1673
rect 1942 1619 1958 1673
rect 1892 1601 1958 1619
rect 1892 1551 1908 1601
rect 1942 1551 1958 1601
rect 1892 1529 1958 1551
rect 1892 1483 1908 1529
rect 1942 1483 1958 1529
rect 1892 1457 1958 1483
rect 1892 1415 1908 1457
rect 1942 1415 1958 1457
rect 1892 1385 1958 1415
rect 1892 1347 1908 1385
rect 1942 1347 1958 1385
rect 1892 1313 1958 1347
rect 1892 1279 1908 1313
rect 1942 1279 1958 1313
rect 1892 1245 1958 1279
rect 1892 1207 1908 1245
rect 1942 1207 1958 1245
rect 1892 1177 1958 1207
rect 1892 1135 1908 1177
rect 1942 1135 1958 1177
rect 1892 1109 1958 1135
rect 1892 1063 1908 1109
rect 1942 1063 1958 1109
rect 1892 1041 1958 1063
rect 1892 991 1908 1041
rect 1942 991 1958 1041
rect 1892 973 1958 991
rect 1892 919 1908 973
rect 1942 919 1958 973
rect 1892 905 1958 919
rect 1892 847 1908 905
rect 1942 847 1958 905
rect 1892 837 1958 847
rect 1892 775 1908 837
rect 1942 775 1958 837
rect 1892 769 1958 775
rect 1892 703 1908 769
rect 1942 703 1958 769
rect 1892 701 1958 703
rect 1892 667 1908 701
rect 1942 667 1958 701
rect 1892 665 1958 667
rect 1892 599 1908 665
rect 1942 599 1958 665
rect 1892 593 1958 599
rect 1892 531 1908 593
rect 1942 531 1958 593
rect 1892 521 1958 531
rect 1892 463 1908 521
rect 1942 463 1958 521
rect 1892 449 1958 463
rect 1892 395 1908 449
rect 1942 395 1958 449
rect 1892 377 1958 395
rect 1892 327 1908 377
rect 1942 327 1958 377
rect 1892 305 1958 327
rect 34 233 100 259
rect 34 191 50 233
rect 84 191 100 233
rect 34 161 100 191
rect 34 123 50 161
rect 84 123 100 161
rect 34 100 100 123
rect 1892 259 1908 305
rect 1942 259 1958 305
rect 1892 233 1958 259
rect 1892 191 1908 233
rect 1942 191 1958 233
rect 1892 161 1958 191
rect 1892 123 1908 161
rect 1942 123 1958 161
rect 1892 100 1958 123
rect 34 84 1958 100
rect 34 50 50 84
rect 84 50 129 84
rect 185 50 197 84
rect 257 50 265 84
rect 329 50 333 84
rect 435 50 439 84
rect 503 50 511 84
rect 571 50 583 84
rect 639 50 655 84
rect 707 50 727 84
rect 775 50 799 84
rect 843 50 871 84
rect 911 50 943 84
rect 979 50 1013 84
rect 1049 50 1081 84
rect 1121 50 1149 84
rect 1193 50 1217 84
rect 1265 50 1285 84
rect 1337 50 1353 84
rect 1409 50 1421 84
rect 1481 50 1489 84
rect 1553 50 1557 84
rect 1659 50 1663 84
rect 1727 50 1735 84
rect 1795 50 1807 84
rect 1863 50 1908 84
rect 1942 50 1958 84
rect 34 34 1958 50
<< viali >>
rect 50 2508 84 2542
rect 151 2508 163 2542
rect 163 2508 185 2542
rect 223 2508 231 2542
rect 231 2508 257 2542
rect 295 2508 299 2542
rect 299 2508 329 2542
rect 367 2508 401 2542
rect 439 2508 469 2542
rect 469 2508 473 2542
rect 511 2508 537 2542
rect 537 2508 545 2542
rect 583 2508 605 2542
rect 605 2508 617 2542
rect 655 2508 673 2542
rect 673 2508 689 2542
rect 727 2508 741 2542
rect 741 2508 761 2542
rect 799 2508 809 2542
rect 809 2508 833 2542
rect 871 2508 877 2542
rect 877 2508 905 2542
rect 943 2508 945 2542
rect 945 2508 977 2542
rect 1015 2508 1047 2542
rect 1047 2508 1049 2542
rect 1087 2508 1115 2542
rect 1115 2508 1121 2542
rect 1159 2508 1183 2542
rect 1183 2508 1193 2542
rect 1231 2508 1251 2542
rect 1251 2508 1265 2542
rect 1303 2508 1319 2542
rect 1319 2508 1337 2542
rect 1375 2508 1387 2542
rect 1387 2508 1409 2542
rect 1447 2508 1455 2542
rect 1455 2508 1481 2542
rect 1519 2508 1523 2542
rect 1523 2508 1553 2542
rect 1591 2508 1625 2542
rect 1663 2508 1693 2542
rect 1693 2508 1697 2542
rect 1735 2508 1761 2542
rect 1761 2508 1769 2542
rect 1807 2508 1829 2542
rect 1829 2508 1841 2542
rect 1908 2508 1942 2542
rect 50 2435 84 2465
rect 50 2431 84 2435
rect 50 2367 84 2393
rect 50 2359 84 2367
rect 50 2299 84 2321
rect 50 2287 84 2299
rect 1908 2435 1942 2465
rect 1908 2431 1942 2435
rect 1908 2367 1942 2393
rect 1908 2359 1942 2367
rect 50 2231 84 2249
rect 50 2215 84 2231
rect 50 2163 84 2177
rect 50 2143 84 2163
rect 50 2095 84 2105
rect 50 2071 84 2095
rect 50 2027 84 2033
rect 50 1999 84 2027
rect 50 1959 84 1961
rect 50 1927 84 1959
rect 50 1857 84 1889
rect 50 1855 84 1857
rect 50 1789 84 1817
rect 50 1783 84 1789
rect 50 1721 84 1745
rect 50 1711 84 1721
rect 50 1653 84 1673
rect 50 1639 84 1653
rect 50 1585 84 1601
rect 50 1567 84 1585
rect 50 1517 84 1529
rect 50 1495 84 1517
rect 50 1449 84 1457
rect 50 1423 84 1449
rect 50 1381 84 1385
rect 50 1351 84 1381
rect 50 1279 84 1313
rect 50 1211 84 1241
rect 50 1207 84 1211
rect 50 1143 84 1169
rect 50 1135 84 1143
rect 50 1075 84 1097
rect 50 1063 84 1075
rect 50 1007 84 1025
rect 50 991 84 1007
rect 50 939 84 953
rect 50 919 84 939
rect 50 871 84 881
rect 50 847 84 871
rect 50 803 84 809
rect 50 775 84 803
rect 50 735 84 737
rect 50 703 84 735
rect 50 633 84 665
rect 50 631 84 633
rect 50 565 84 593
rect 50 559 84 565
rect 50 497 84 521
rect 50 487 84 497
rect 50 429 84 449
rect 50 415 84 429
rect 50 361 84 377
rect 50 343 84 361
rect 50 293 84 305
rect 50 271 84 293
rect 276 2282 310 2316
rect 367 2282 401 2316
rect 439 2282 469 2316
rect 469 2282 473 2316
rect 511 2282 537 2316
rect 537 2282 545 2316
rect 583 2282 605 2316
rect 605 2282 617 2316
rect 655 2282 673 2316
rect 673 2282 689 2316
rect 727 2282 741 2316
rect 741 2282 761 2316
rect 799 2282 809 2316
rect 809 2282 833 2316
rect 871 2282 877 2316
rect 877 2282 905 2316
rect 943 2282 945 2316
rect 945 2282 977 2316
rect 1015 2282 1047 2316
rect 1047 2282 1049 2316
rect 1087 2282 1115 2316
rect 1115 2282 1121 2316
rect 1159 2282 1183 2316
rect 1183 2282 1193 2316
rect 1231 2282 1251 2316
rect 1251 2282 1265 2316
rect 1303 2282 1319 2316
rect 1319 2282 1337 2316
rect 1375 2282 1387 2316
rect 1387 2282 1409 2316
rect 1447 2282 1455 2316
rect 1455 2282 1481 2316
rect 1519 2282 1523 2316
rect 1523 2282 1553 2316
rect 1591 2282 1625 2316
rect 1682 2282 1716 2316
rect 276 2197 310 2213
rect 276 2179 310 2197
rect 276 2129 310 2141
rect 276 2107 310 2129
rect 276 2061 310 2069
rect 276 2035 310 2061
rect 276 1993 310 1997
rect 276 1963 310 1993
rect 276 1891 310 1925
rect 1682 2197 1716 2213
rect 1682 2179 1716 2197
rect 1682 2129 1716 2141
rect 1682 2107 1716 2129
rect 1682 2061 1716 2069
rect 1682 2035 1716 2061
rect 1682 1993 1716 1997
rect 1682 1963 1716 1993
rect 276 1823 310 1853
rect 276 1819 310 1823
rect 276 1755 310 1781
rect 276 1747 310 1755
rect 276 1687 310 1709
rect 276 1675 310 1687
rect 276 1619 310 1637
rect 276 1603 310 1619
rect 276 1551 310 1565
rect 276 1531 310 1551
rect 276 1483 310 1493
rect 276 1459 310 1483
rect 276 1415 310 1421
rect 276 1387 310 1415
rect 276 1347 310 1349
rect 276 1315 310 1347
rect 276 1245 310 1277
rect 276 1243 310 1245
rect 276 1177 310 1205
rect 276 1171 310 1177
rect 276 1109 310 1133
rect 276 1099 310 1109
rect 276 1041 310 1061
rect 276 1027 310 1041
rect 276 973 310 989
rect 276 955 310 973
rect 276 905 310 917
rect 276 883 310 905
rect 276 837 310 845
rect 276 811 310 837
rect 276 769 310 773
rect 276 739 310 769
rect 276 667 310 701
rect 678 1880 712 1914
rect 763 1880 775 1914
rect 775 1880 797 1914
rect 835 1880 843 1914
rect 843 1880 869 1914
rect 907 1880 911 1914
rect 911 1880 941 1914
rect 979 1880 1013 1914
rect 1051 1880 1081 1914
rect 1081 1880 1085 1914
rect 1123 1880 1149 1914
rect 1149 1880 1157 1914
rect 1195 1880 1217 1914
rect 1217 1880 1229 1914
rect 1280 1880 1314 1914
rect 678 1789 712 1817
rect 678 1783 712 1789
rect 678 1721 712 1745
rect 678 1711 712 1721
rect 1280 1789 1314 1817
rect 1280 1783 1314 1789
rect 1280 1721 1314 1745
rect 1280 1711 1314 1721
rect 678 1653 712 1673
rect 678 1639 712 1653
rect 678 1585 712 1601
rect 678 1567 712 1585
rect 678 1517 712 1529
rect 678 1495 712 1517
rect 678 1449 712 1457
rect 678 1423 712 1449
rect 678 1381 712 1385
rect 678 1351 712 1381
rect 678 1279 712 1313
rect 678 1211 712 1241
rect 678 1207 712 1211
rect 678 1143 712 1169
rect 678 1135 712 1143
rect 678 1075 712 1097
rect 678 1063 712 1075
rect 678 1007 712 1025
rect 678 991 712 1007
rect 678 939 712 953
rect 678 919 712 939
rect 907 1653 1085 1673
rect 907 939 911 1653
rect 911 939 1081 1653
rect 1081 939 1085 1653
rect 907 919 1085 939
rect 1280 1653 1314 1673
rect 1280 1639 1314 1653
rect 1280 1585 1314 1601
rect 1280 1567 1314 1585
rect 1280 1517 1314 1529
rect 1280 1495 1314 1517
rect 1280 1449 1314 1457
rect 1280 1423 1314 1449
rect 1280 1381 1314 1385
rect 1280 1351 1314 1381
rect 1280 1279 1314 1313
rect 1280 1211 1314 1241
rect 1280 1207 1314 1211
rect 1280 1143 1314 1169
rect 1280 1135 1314 1143
rect 1280 1075 1314 1097
rect 1280 1063 1314 1075
rect 1280 1007 1314 1025
rect 1280 991 1314 1007
rect 1280 939 1314 953
rect 1280 919 1314 939
rect 678 871 712 881
rect 678 847 712 871
rect 678 803 712 809
rect 678 775 712 803
rect 1280 871 1314 881
rect 1280 847 1314 871
rect 1280 803 1314 809
rect 1280 775 1314 803
rect 678 678 712 712
rect 763 678 775 712
rect 775 678 797 712
rect 835 678 843 712
rect 843 678 869 712
rect 907 678 911 712
rect 911 678 941 712
rect 979 678 1013 712
rect 1051 678 1081 712
rect 1081 678 1085 712
rect 1123 678 1149 712
rect 1149 678 1157 712
rect 1195 678 1217 712
rect 1217 678 1229 712
rect 1280 678 1314 712
rect 1682 1891 1716 1925
rect 1682 1823 1716 1853
rect 1682 1819 1716 1823
rect 1682 1755 1716 1781
rect 1682 1747 1716 1755
rect 1682 1687 1716 1709
rect 1682 1675 1716 1687
rect 1682 1619 1716 1637
rect 1682 1603 1716 1619
rect 1682 1551 1716 1565
rect 1682 1531 1716 1551
rect 1682 1483 1716 1493
rect 1682 1459 1716 1483
rect 1682 1415 1716 1421
rect 1682 1387 1716 1415
rect 1682 1347 1716 1349
rect 1682 1315 1716 1347
rect 1682 1245 1716 1277
rect 1682 1243 1716 1245
rect 1682 1177 1716 1205
rect 1682 1171 1716 1177
rect 1682 1109 1716 1133
rect 1682 1099 1716 1109
rect 1682 1041 1716 1061
rect 1682 1027 1716 1041
rect 1682 973 1716 989
rect 1682 955 1716 973
rect 1682 905 1716 917
rect 1682 883 1716 905
rect 1682 837 1716 845
rect 1682 811 1716 837
rect 1682 769 1716 773
rect 1682 739 1716 769
rect 276 599 310 629
rect 276 595 310 599
rect 276 531 310 557
rect 276 523 310 531
rect 276 463 310 485
rect 276 451 310 463
rect 276 395 310 413
rect 276 379 310 395
rect 1682 667 1716 701
rect 1682 599 1716 629
rect 1682 595 1716 599
rect 1682 531 1716 557
rect 1682 523 1716 531
rect 1682 463 1716 485
rect 1682 451 1716 463
rect 1682 395 1716 413
rect 1682 379 1716 395
rect 276 276 310 310
rect 367 276 401 310
rect 439 276 469 310
rect 469 276 473 310
rect 511 276 537 310
rect 537 276 545 310
rect 583 276 605 310
rect 605 276 617 310
rect 655 276 673 310
rect 673 276 689 310
rect 727 276 741 310
rect 741 276 761 310
rect 799 276 809 310
rect 809 276 833 310
rect 871 276 877 310
rect 877 276 905 310
rect 943 276 945 310
rect 945 276 977 310
rect 1015 276 1047 310
rect 1047 276 1049 310
rect 1087 276 1115 310
rect 1115 276 1121 310
rect 1159 276 1183 310
rect 1183 276 1193 310
rect 1231 276 1251 310
rect 1251 276 1265 310
rect 1303 276 1319 310
rect 1319 276 1337 310
rect 1375 276 1387 310
rect 1387 276 1409 310
rect 1447 276 1455 310
rect 1455 276 1481 310
rect 1519 276 1523 310
rect 1523 276 1553 310
rect 1591 276 1625 310
rect 1682 276 1716 310
rect 1908 2299 1942 2321
rect 1908 2287 1942 2299
rect 1908 2231 1942 2249
rect 1908 2215 1942 2231
rect 1908 2163 1942 2177
rect 1908 2143 1942 2163
rect 1908 2095 1942 2105
rect 1908 2071 1942 2095
rect 1908 2027 1942 2033
rect 1908 1999 1942 2027
rect 1908 1959 1942 1961
rect 1908 1927 1942 1959
rect 1908 1857 1942 1889
rect 1908 1855 1942 1857
rect 1908 1789 1942 1817
rect 1908 1783 1942 1789
rect 1908 1721 1942 1745
rect 1908 1711 1942 1721
rect 1908 1653 1942 1673
rect 1908 1639 1942 1653
rect 1908 1585 1942 1601
rect 1908 1567 1942 1585
rect 1908 1517 1942 1529
rect 1908 1495 1942 1517
rect 1908 1449 1942 1457
rect 1908 1423 1942 1449
rect 1908 1381 1942 1385
rect 1908 1351 1942 1381
rect 1908 1279 1942 1313
rect 1908 1211 1942 1241
rect 1908 1207 1942 1211
rect 1908 1143 1942 1169
rect 1908 1135 1942 1143
rect 1908 1075 1942 1097
rect 1908 1063 1942 1075
rect 1908 1007 1942 1025
rect 1908 991 1942 1007
rect 1908 939 1942 953
rect 1908 919 1942 939
rect 1908 871 1942 881
rect 1908 847 1942 871
rect 1908 803 1942 809
rect 1908 775 1942 803
rect 1908 735 1942 737
rect 1908 703 1942 735
rect 1908 633 1942 665
rect 1908 631 1942 633
rect 1908 565 1942 593
rect 1908 559 1942 565
rect 1908 497 1942 521
rect 1908 487 1942 497
rect 1908 429 1942 449
rect 1908 415 1942 429
rect 1908 361 1942 377
rect 1908 343 1942 361
rect 50 225 84 233
rect 50 199 84 225
rect 50 157 84 161
rect 50 127 84 157
rect 1908 293 1942 305
rect 1908 271 1942 293
rect 1908 225 1942 233
rect 1908 199 1942 225
rect 1908 157 1942 161
rect 1908 127 1942 157
rect 50 50 84 84
rect 151 50 163 84
rect 163 50 185 84
rect 223 50 231 84
rect 231 50 257 84
rect 295 50 299 84
rect 299 50 329 84
rect 367 50 401 84
rect 439 50 469 84
rect 469 50 473 84
rect 511 50 537 84
rect 537 50 545 84
rect 583 50 605 84
rect 605 50 617 84
rect 655 50 673 84
rect 673 50 689 84
rect 727 50 741 84
rect 741 50 761 84
rect 799 50 809 84
rect 809 50 833 84
rect 871 50 877 84
rect 877 50 905 84
rect 943 50 945 84
rect 945 50 977 84
rect 1015 50 1047 84
rect 1047 50 1049 84
rect 1087 50 1115 84
rect 1115 50 1121 84
rect 1159 50 1183 84
rect 1183 50 1193 84
rect 1231 50 1251 84
rect 1251 50 1265 84
rect 1303 50 1319 84
rect 1319 50 1337 84
rect 1375 50 1387 84
rect 1387 50 1409 84
rect 1447 50 1455 84
rect 1455 50 1481 84
rect 1519 50 1523 84
rect 1523 50 1553 84
rect 1591 50 1625 84
rect 1663 50 1693 84
rect 1693 50 1697 84
rect 1735 50 1761 84
rect 1761 50 1769 84
rect 1807 50 1829 84
rect 1829 50 1841 84
rect 1908 50 1942 84
<< metal1 >>
rect 38 2542 1954 2554
rect 38 2508 50 2542
rect 84 2508 151 2542
rect 185 2508 223 2542
rect 257 2508 295 2542
rect 329 2508 367 2542
rect 401 2508 439 2542
rect 473 2508 511 2542
rect 545 2508 583 2542
rect 617 2508 655 2542
rect 689 2508 727 2542
rect 761 2508 799 2542
rect 833 2508 871 2542
rect 905 2508 943 2542
rect 977 2508 1015 2542
rect 1049 2508 1087 2542
rect 1121 2508 1159 2542
rect 1193 2508 1231 2542
rect 1265 2508 1303 2542
rect 1337 2508 1375 2542
rect 1409 2508 1447 2542
rect 1481 2508 1519 2542
rect 1553 2508 1591 2542
rect 1625 2508 1663 2542
rect 1697 2508 1735 2542
rect 1769 2508 1807 2542
rect 1841 2508 1908 2542
rect 1942 2508 1954 2542
rect 38 2496 1954 2508
rect 38 2465 96 2496
rect 38 2431 50 2465
rect 84 2431 96 2465
rect 38 2393 96 2431
rect 38 2359 50 2393
rect 84 2359 96 2393
rect 38 2321 96 2359
rect 1896 2465 1954 2496
rect 1896 2431 1908 2465
rect 1942 2431 1954 2465
rect 1896 2393 1954 2431
rect 1896 2359 1908 2393
rect 1942 2359 1954 2393
rect 38 2287 50 2321
rect 84 2287 96 2321
rect 38 2249 96 2287
rect 38 2215 50 2249
rect 84 2215 96 2249
rect 38 2177 96 2215
rect 38 2143 50 2177
rect 84 2143 96 2177
rect 38 2105 96 2143
rect 38 2071 50 2105
rect 84 2071 96 2105
rect 38 2033 96 2071
rect 38 1999 50 2033
rect 84 1999 96 2033
rect 38 1961 96 1999
rect 38 1927 50 1961
rect 84 1927 96 1961
rect 38 1889 96 1927
rect 38 1855 50 1889
rect 84 1855 96 1889
rect 38 1817 96 1855
rect 38 1783 50 1817
rect 84 1783 96 1817
rect 38 1745 96 1783
rect 38 1711 50 1745
rect 84 1711 96 1745
rect 38 1673 96 1711
rect 38 1639 50 1673
rect 84 1639 96 1673
rect 38 1601 96 1639
rect 38 1567 50 1601
rect 84 1567 96 1601
rect 38 1529 96 1567
rect 38 1495 50 1529
rect 84 1495 96 1529
rect 38 1457 96 1495
rect 38 1423 50 1457
rect 84 1423 96 1457
rect 38 1385 96 1423
rect 38 1351 50 1385
rect 84 1351 96 1385
rect 38 1313 96 1351
rect 38 1279 50 1313
rect 84 1279 96 1313
rect 38 1241 96 1279
rect 38 1207 50 1241
rect 84 1207 96 1241
rect 38 1169 96 1207
rect 38 1135 50 1169
rect 84 1135 96 1169
rect 38 1097 96 1135
rect 38 1063 50 1097
rect 84 1063 96 1097
rect 38 1025 96 1063
rect 38 991 50 1025
rect 84 991 96 1025
rect 38 953 96 991
rect 38 919 50 953
rect 84 919 96 953
rect 38 881 96 919
rect 38 847 50 881
rect 84 847 96 881
rect 38 809 96 847
rect 38 775 50 809
rect 84 775 96 809
rect 38 737 96 775
rect 38 703 50 737
rect 84 703 96 737
rect 38 665 96 703
rect 38 631 50 665
rect 84 631 96 665
rect 38 593 96 631
rect 38 559 50 593
rect 84 559 96 593
rect 38 521 96 559
rect 38 487 50 521
rect 84 487 96 521
rect 38 449 96 487
rect 38 415 50 449
rect 84 415 96 449
rect 38 377 96 415
rect 38 343 50 377
rect 84 343 96 377
rect 38 305 96 343
rect 38 271 50 305
rect 84 271 96 305
rect 38 233 96 271
rect 264 2316 1728 2328
rect 264 2282 276 2316
rect 310 2282 367 2316
rect 401 2282 439 2316
rect 473 2282 511 2316
rect 545 2282 583 2316
rect 617 2282 655 2316
rect 689 2282 727 2316
rect 761 2282 799 2316
rect 833 2282 871 2316
rect 905 2282 943 2316
rect 977 2282 1015 2316
rect 1049 2282 1087 2316
rect 1121 2282 1159 2316
rect 1193 2282 1231 2316
rect 1265 2282 1303 2316
rect 1337 2282 1375 2316
rect 1409 2282 1447 2316
rect 1481 2282 1519 2316
rect 1553 2282 1591 2316
rect 1625 2282 1682 2316
rect 1716 2282 1728 2316
rect 264 2270 1728 2282
rect 264 2213 322 2270
rect 264 2179 276 2213
rect 310 2179 322 2213
rect 264 2141 322 2179
rect 264 2107 276 2141
rect 310 2107 322 2141
rect 264 2069 322 2107
rect 264 2035 276 2069
rect 310 2035 322 2069
rect 264 1997 322 2035
rect 264 1963 276 1997
rect 310 1963 322 1997
rect 264 1925 322 1963
rect 1670 2213 1728 2270
rect 1670 2179 1682 2213
rect 1716 2179 1728 2213
rect 1670 2141 1728 2179
rect 1670 2107 1682 2141
rect 1716 2107 1728 2141
rect 1670 2069 1728 2107
rect 1670 2035 1682 2069
rect 1716 2035 1728 2069
rect 1670 1997 1728 2035
rect 1670 1963 1682 1997
rect 1716 1963 1728 1997
rect 264 1891 276 1925
rect 310 1891 322 1925
rect 264 1853 322 1891
rect 264 1819 276 1853
rect 310 1819 322 1853
rect 264 1781 322 1819
rect 264 1747 276 1781
rect 310 1747 322 1781
rect 264 1709 322 1747
rect 264 1675 276 1709
rect 310 1675 322 1709
rect 264 1637 322 1675
rect 264 1603 276 1637
rect 310 1603 322 1637
rect 264 1565 322 1603
rect 264 1531 276 1565
rect 310 1531 322 1565
rect 264 1493 322 1531
rect 264 1459 276 1493
rect 310 1459 322 1493
rect 264 1421 322 1459
rect 264 1387 276 1421
rect 310 1387 322 1421
rect 264 1349 322 1387
rect 264 1315 276 1349
rect 310 1315 322 1349
rect 264 1277 322 1315
rect 264 1243 276 1277
rect 310 1243 322 1277
rect 264 1205 322 1243
rect 264 1171 276 1205
rect 310 1171 322 1205
rect 264 1133 322 1171
rect 264 1099 276 1133
rect 310 1099 322 1133
rect 264 1061 322 1099
rect 264 1027 276 1061
rect 310 1027 322 1061
rect 264 989 322 1027
rect 264 955 276 989
rect 310 955 322 989
rect 264 917 322 955
rect 264 883 276 917
rect 310 883 322 917
rect 264 845 322 883
rect 264 811 276 845
rect 310 811 322 845
rect 264 773 322 811
rect 264 739 276 773
rect 310 739 322 773
rect 264 701 322 739
rect 264 667 276 701
rect 310 667 322 701
rect 264 629 322 667
rect 666 1914 1326 1926
rect 666 1880 678 1914
rect 712 1880 763 1914
rect 797 1880 835 1914
rect 869 1880 907 1914
rect 941 1880 979 1914
rect 1013 1880 1051 1914
rect 1085 1880 1123 1914
rect 1157 1880 1195 1914
rect 1229 1880 1280 1914
rect 1314 1880 1326 1914
rect 666 1868 1326 1880
rect 666 1817 724 1868
rect 666 1783 678 1817
rect 712 1783 724 1817
rect 666 1745 724 1783
rect 666 1711 678 1745
rect 712 1711 724 1745
rect 666 1673 724 1711
rect 1268 1817 1326 1868
rect 1268 1783 1280 1817
rect 1314 1783 1326 1817
rect 1268 1745 1326 1783
rect 1268 1711 1280 1745
rect 1314 1711 1326 1745
rect 666 1639 678 1673
rect 712 1639 724 1673
rect 666 1601 724 1639
rect 666 1567 678 1601
rect 712 1567 724 1601
rect 666 1529 724 1567
rect 666 1495 678 1529
rect 712 1495 724 1529
rect 666 1457 724 1495
rect 666 1423 678 1457
rect 712 1423 724 1457
rect 666 1385 724 1423
rect 666 1351 678 1385
rect 712 1351 724 1385
rect 666 1313 724 1351
rect 666 1279 678 1313
rect 712 1279 724 1313
rect 666 1241 724 1279
rect 666 1207 678 1241
rect 712 1207 724 1241
rect 666 1169 724 1207
rect 666 1135 678 1169
rect 712 1135 724 1169
rect 666 1097 724 1135
rect 666 1063 678 1097
rect 712 1063 724 1097
rect 666 1025 724 1063
rect 666 991 678 1025
rect 712 991 724 1025
rect 666 953 724 991
rect 666 919 678 953
rect 712 919 724 953
rect 666 881 724 919
rect 895 1673 1097 1685
rect 895 919 907 1673
rect 1085 919 1097 1673
rect 895 907 1097 919
rect 1268 1673 1326 1711
rect 1268 1639 1280 1673
rect 1314 1639 1326 1673
rect 1268 1601 1326 1639
rect 1268 1567 1280 1601
rect 1314 1567 1326 1601
rect 1268 1529 1326 1567
rect 1268 1495 1280 1529
rect 1314 1495 1326 1529
rect 1268 1457 1326 1495
rect 1268 1423 1280 1457
rect 1314 1423 1326 1457
rect 1268 1385 1326 1423
rect 1268 1351 1280 1385
rect 1314 1351 1326 1385
rect 1268 1313 1326 1351
rect 1268 1279 1280 1313
rect 1314 1279 1326 1313
rect 1268 1241 1326 1279
rect 1268 1207 1280 1241
rect 1314 1207 1326 1241
rect 1268 1169 1326 1207
rect 1268 1135 1280 1169
rect 1314 1135 1326 1169
rect 1268 1097 1326 1135
rect 1268 1063 1280 1097
rect 1314 1063 1326 1097
rect 1268 1025 1326 1063
rect 1268 991 1280 1025
rect 1314 991 1326 1025
rect 1268 953 1326 991
rect 1268 919 1280 953
rect 1314 919 1326 953
rect 666 847 678 881
rect 712 847 724 881
rect 666 809 724 847
rect 666 775 678 809
rect 712 775 724 809
rect 666 724 724 775
rect 1268 881 1326 919
rect 1268 847 1280 881
rect 1314 847 1326 881
rect 1268 809 1326 847
rect 1268 775 1280 809
rect 1314 775 1326 809
rect 1268 724 1326 775
rect 666 712 1326 724
rect 666 678 678 712
rect 712 678 763 712
rect 797 678 835 712
rect 869 678 907 712
rect 941 678 979 712
rect 1013 678 1051 712
rect 1085 678 1123 712
rect 1157 678 1195 712
rect 1229 678 1280 712
rect 1314 678 1326 712
rect 666 666 1326 678
rect 1670 1925 1728 1963
rect 1670 1891 1682 1925
rect 1716 1891 1728 1925
rect 1670 1853 1728 1891
rect 1670 1819 1682 1853
rect 1716 1819 1728 1853
rect 1670 1781 1728 1819
rect 1670 1747 1682 1781
rect 1716 1747 1728 1781
rect 1670 1709 1728 1747
rect 1670 1675 1682 1709
rect 1716 1675 1728 1709
rect 1670 1637 1728 1675
rect 1670 1603 1682 1637
rect 1716 1603 1728 1637
rect 1670 1565 1728 1603
rect 1670 1531 1682 1565
rect 1716 1531 1728 1565
rect 1670 1493 1728 1531
rect 1670 1459 1682 1493
rect 1716 1459 1728 1493
rect 1670 1421 1728 1459
rect 1670 1387 1682 1421
rect 1716 1387 1728 1421
rect 1670 1349 1728 1387
rect 1670 1315 1682 1349
rect 1716 1315 1728 1349
rect 1670 1277 1728 1315
rect 1670 1243 1682 1277
rect 1716 1243 1728 1277
rect 1670 1205 1728 1243
rect 1670 1171 1682 1205
rect 1716 1171 1728 1205
rect 1670 1133 1728 1171
rect 1670 1099 1682 1133
rect 1716 1099 1728 1133
rect 1670 1061 1728 1099
rect 1670 1027 1682 1061
rect 1716 1027 1728 1061
rect 1670 989 1728 1027
rect 1670 955 1682 989
rect 1716 955 1728 989
rect 1670 917 1728 955
rect 1670 883 1682 917
rect 1716 883 1728 917
rect 1670 845 1728 883
rect 1670 811 1682 845
rect 1716 811 1728 845
rect 1670 773 1728 811
rect 1670 739 1682 773
rect 1716 739 1728 773
rect 1670 701 1728 739
rect 1670 667 1682 701
rect 1716 667 1728 701
rect 264 595 276 629
rect 310 595 322 629
rect 264 557 322 595
rect 264 523 276 557
rect 310 523 322 557
rect 264 485 322 523
rect 264 451 276 485
rect 310 451 322 485
rect 264 413 322 451
rect 264 379 276 413
rect 310 379 322 413
rect 264 322 322 379
rect 1670 629 1728 667
rect 1670 595 1682 629
rect 1716 595 1728 629
rect 1670 557 1728 595
rect 1670 523 1682 557
rect 1716 523 1728 557
rect 1670 485 1728 523
rect 1670 451 1682 485
rect 1716 451 1728 485
rect 1670 413 1728 451
rect 1670 379 1682 413
rect 1716 379 1728 413
rect 1670 322 1728 379
rect 264 310 1728 322
rect 264 276 276 310
rect 310 276 367 310
rect 401 276 439 310
rect 473 276 511 310
rect 545 276 583 310
rect 617 276 655 310
rect 689 276 727 310
rect 761 276 799 310
rect 833 276 871 310
rect 905 276 943 310
rect 977 276 1015 310
rect 1049 276 1087 310
rect 1121 276 1159 310
rect 1193 276 1231 310
rect 1265 276 1303 310
rect 1337 276 1375 310
rect 1409 276 1447 310
rect 1481 276 1519 310
rect 1553 276 1591 310
rect 1625 276 1682 310
rect 1716 276 1728 310
rect 264 264 1728 276
rect 1896 2321 1954 2359
rect 1896 2287 1908 2321
rect 1942 2287 1954 2321
rect 1896 2249 1954 2287
rect 1896 2215 1908 2249
rect 1942 2215 1954 2249
rect 1896 2177 1954 2215
rect 1896 2143 1908 2177
rect 1942 2143 1954 2177
rect 1896 2105 1954 2143
rect 1896 2071 1908 2105
rect 1942 2071 1954 2105
rect 1896 2033 1954 2071
rect 1896 1999 1908 2033
rect 1942 1999 1954 2033
rect 1896 1961 1954 1999
rect 1896 1927 1908 1961
rect 1942 1927 1954 1961
rect 1896 1889 1954 1927
rect 1896 1855 1908 1889
rect 1942 1855 1954 1889
rect 1896 1817 1954 1855
rect 1896 1783 1908 1817
rect 1942 1783 1954 1817
rect 1896 1745 1954 1783
rect 1896 1711 1908 1745
rect 1942 1711 1954 1745
rect 1896 1673 1954 1711
rect 1896 1639 1908 1673
rect 1942 1639 1954 1673
rect 1896 1601 1954 1639
rect 1896 1567 1908 1601
rect 1942 1567 1954 1601
rect 1896 1529 1954 1567
rect 1896 1495 1908 1529
rect 1942 1495 1954 1529
rect 1896 1457 1954 1495
rect 1896 1423 1908 1457
rect 1942 1423 1954 1457
rect 1896 1385 1954 1423
rect 1896 1351 1908 1385
rect 1942 1351 1954 1385
rect 1896 1313 1954 1351
rect 1896 1279 1908 1313
rect 1942 1279 1954 1313
rect 1896 1241 1954 1279
rect 1896 1207 1908 1241
rect 1942 1207 1954 1241
rect 1896 1169 1954 1207
rect 1896 1135 1908 1169
rect 1942 1135 1954 1169
rect 1896 1097 1954 1135
rect 1896 1063 1908 1097
rect 1942 1063 1954 1097
rect 1896 1025 1954 1063
rect 1896 991 1908 1025
rect 1942 991 1954 1025
rect 1896 953 1954 991
rect 1896 919 1908 953
rect 1942 919 1954 953
rect 1896 881 1954 919
rect 1896 847 1908 881
rect 1942 847 1954 881
rect 1896 809 1954 847
rect 1896 775 1908 809
rect 1942 775 1954 809
rect 1896 737 1954 775
rect 1896 703 1908 737
rect 1942 703 1954 737
rect 1896 665 1954 703
rect 1896 631 1908 665
rect 1942 631 1954 665
rect 1896 593 1954 631
rect 1896 559 1908 593
rect 1942 559 1954 593
rect 1896 521 1954 559
rect 1896 487 1908 521
rect 1942 487 1954 521
rect 1896 449 1954 487
rect 1896 415 1908 449
rect 1942 415 1954 449
rect 1896 377 1954 415
rect 1896 343 1908 377
rect 1942 343 1954 377
rect 1896 305 1954 343
rect 1896 271 1908 305
rect 1942 271 1954 305
rect 38 199 50 233
rect 84 199 96 233
rect 38 161 96 199
rect 38 127 50 161
rect 84 127 96 161
rect 38 96 96 127
rect 1896 233 1954 271
rect 1896 199 1908 233
rect 1942 199 1954 233
rect 1896 161 1954 199
rect 1896 127 1908 161
rect 1942 127 1954 161
rect 1896 96 1954 127
rect 38 84 1954 96
rect 38 50 50 84
rect 84 50 151 84
rect 185 50 223 84
rect 257 50 295 84
rect 329 50 367 84
rect 401 50 439 84
rect 473 50 511 84
rect 545 50 583 84
rect 617 50 655 84
rect 689 50 727 84
rect 761 50 799 84
rect 833 50 871 84
rect 905 50 943 84
rect 977 50 1015 84
rect 1049 50 1087 84
rect 1121 50 1159 84
rect 1193 50 1231 84
rect 1265 50 1303 84
rect 1337 50 1375 84
rect 1409 50 1447 84
rect 1481 50 1519 84
rect 1553 50 1591 84
rect 1625 50 1663 84
rect 1697 50 1735 84
rect 1769 50 1807 84
rect 1841 50 1908 84
rect 1942 50 1954 84
rect 38 38 1954 50
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 8888328
string GDS_START 8840764
string path 7.850 12.350 7.850 56.950 41.950 56.950 41.950 7.850 3.350 7.850 
<< end >>
